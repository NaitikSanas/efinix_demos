
//
// Verific Verilog Description of module mipi_pi_top
//

module mipi_pi_top (i_arstn, mipi_pclk, mipi_inst1_DPHY_RSTN, mipi_inst1_RSTN, 
            mipi_inst1_VC_ENA, mipi_inst1_LANES, mipi_inst1_CLEAR, mipi_inst1_HSYNC, 
            mipi_inst1_VSYNC, mipi_inst1_CNT, mipi_inst1_VALID, mipi_inst1_TYPE, 
            mipi_inst1_DATA, mipi_inst1_VC, mipi_inst1_ERR, mipi_inst2_DPHY_RSTN, 
            mipi_inst2_RSTN, mipi_inst2_VALID, mipi_inst2_HSYNC, mipi_inst2_VSYNC, 
            mipi_inst2_DATA, mipi_inst2_TYPE, mipi_inst2_LANES, mipi_inst2_FRAME_MODE, 
            mipi_inst2_HRES, mipi_inst2_VC, mipi_inst2_ULPS_ENTER, mipi_inst2_ULPS_EXIT, 
            mipi_inst2_ULPS_CLK_ENTER, mipi_inst2_ULPS_CLK_EXIT, sys_clk, 
            rx_status, standby, rx_status2, rx_status3, key1, key2);
    input i_arstn /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_pclk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi_inst1_DPHY_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst1_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]mipi_inst1_VC_ENA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]mipi_inst1_LANES /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst1_CLEAR /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input [3:0]mipi_inst1_HSYNC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_inst1_VSYNC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [3:0]mipi_inst1_CNT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input mipi_inst1_VALID /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [5:0]mipi_inst1_TYPE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [63:0]mipi_inst1_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [1:0]mipi_inst1_VC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input [17:0]mipi_inst1_ERR /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output mipi_inst2_DPHY_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst2_RSTN /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst2_VALID /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst2_HSYNC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst2_VSYNC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [63:0]mipi_inst2_DATA /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [5:0]mipi_inst2_TYPE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]mipi_inst2_LANES /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst2_FRAME_MODE /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [15:0]mipi_inst2_HRES /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [1:0]mipi_inst2_VC /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]mipi_inst2_ULPS_ENTER /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output [3:0]mipi_inst2_ULPS_EXIT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst2_ULPS_CLK_ENTER /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output mipi_inst2_ULPS_CLK_EXIT /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input sys_clk /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    output rx_status /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output standby /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output rx_status2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    output rx_status3 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    input key1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    input key2 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    
    
    wire \r_mipi_rx_data_1P[35] , \r_mipi_rx_data_1P[34] , \r_mipi_rx_data_1P[21] , 
        \r_mipi_rx_data_1P[20] , \r_mipi_rx_data_1P[39] , \r_mipi_rx_data_1P[38] , 
        \r_mipi_rx_data_1P[37] , \r_mipi_rx_data_1P[36] , \r_mipi_rx_data_1P[19] , 
        \r_mipi_rx_data_1P[18] , \r_mipi_rx_data_1P[17] , \r_mipi_rx_data_1P[16] , 
        \r_mipi_rx_data_1P[15] , \r_mipi_rx_data_1P[14] , \r_mipi_rx_data_1P[13] , 
        \r_mipi_rx_data_1P[12] , \r_mipi_rx_data_1P[11] , \r_mipi_rx_data_1P[23] , 
        \r_mipi_rx_data_1P[10] , \r_mipi_rx_data_1P[9] , \r_mipi_rx_data_1P[8] , 
        \r_mipi_rx_data_1P[7] , \r_mipi_rx_data_1P[22] , \r_mipi_rx_data_1P[6] , 
        \r_mipi_rx_data_1P[5] , \r_mipi_rx_data_1P[4] , \r_mipi_rx_data_1P[3] , 
        \r_mipi_rx_data_1P[2] , \r_mipi_rx_data_1P[1] , \r_mipi_rx_data_1P[33] , 
        n141, n142, \r_mipi_rx_data_1P[0] , \r_mipi_rx_data_1P[32] , 
        \r_mipi_rx_data_1P[31] , r_mipi_rx_valid_1P_2, \key1_counter[0]_2 , 
        \r_mipi_rx_data_1P[30] , \r_mipi_rx_data_1P[29] , n150, n151, 
        \r_mipi_rx_data_1P[28] , n153, n154, n155, n156, n157, n158_2, 
        n159_2, n160_2, n161_2, \key2_counter[0] , \r_mipi_rx_data_1P[25] , 
        \r_mipi_rx_data_1P[24] , \red_gain[0] , \r_waddr_1P[0]_2 , n167_2, 
        n168_2, \r_mipi_rx_data_1P[27] , \r_mipi_rx_data_1P[26] , n171_2, 
        n172_2, n173_2, n174_2, n175_2, n176_2, \r_raddr_1P[0]_2 , 
        r_rden_1P_2, n179_2, n180_2, \r_mipi_rx_hsync_1P[0]_2 , \key1_counter[1] , 
        \key1_counter[2] , \key1_counter[3] , \key1_counter[4] , \key1_counter[5] , 
        \key1_counter[6] , \key1_counter[7] , \key1_counter[8] , \key1_counter[9] , 
        \key1_counter[10] , \key1_counter[11] , \key1_counter[12] , \key1_counter[13] , 
        \key1_counter[14] , \key1_counter[15] , n198, n199, n200, 
        n201, n202, n203, n204, n205, n206, n207, n208, n209, 
        n210, n211, n212, n213, n214, n215, n216, n217, n218, 
        n219, n220, n221, n222, n223, n224, n225, n226, n227, 
        n228, n229, n230, n231, n232, n233, n234, n235, n236, 
        n237, n238, n239, n240, n241, n242, n243, n244, n245, 
        n246, n247, n248, n249, n250, n251, n252, n253, n254, 
        n255, n256, n257, n258, n259, n260, n261, n262, n263, 
        n264, n265, n266, n267, n268, n269, n270, n271_2, n272, 
        n273, n274, n275, n276, n277, n278, n279, n280, n281, 
        n282, n283, n284, n285, n286, n287, n288, n289, \key2_counter[1] , 
        \key2_counter[2] , \key2_counter[3] , \key2_counter[4] , \key2_counter[5] , 
        \key2_counter[6] , \key2_counter[7] , \key2_counter[8] , \key2_counter[9] , 
        \key2_counter[10] , \key2_counter[11] , \key2_counter[12] , \key2_counter[13] , 
        \key2_counter[14] , \key2_counter[15] , \red_gain[1] , \red_gain[2] , 
        \green_gain[2] , n308, n309, \r_waddr_1P[1]_2 , \r_waddr_1P[2]_2 , 
        \r_waddr_1P[3]_2 , \r_waddr_1P[4]_2 , \r_waddr_1P[5]_2 , \r_waddr_1P[6]_2 , 
        \r_waddr_1P[7]_2 , \r_waddr_1P[8]_2 , \r_waddr_1P[9]_2 , \r_waddr_1P[10]_2 , 
        \r_waddr_1P[11]_2 , \r_waddr_1P[12]_2 , n322, n323, n324, 
        n325, n326, n327, n328, n329, n330, n331, n332, n333, 
        n334, n335, n336, n337, n338, n339, n340, n341, n342, 
        n343, n344, n345, n346, n347, n348, n349, n350, n351, 
        n352, n353, n354, n355, n356, n357, n358, n359, n360, 
        n361, n362, n363, n364, n365_2, n366_2, n367_2, n368_2, 
        n369_2, n370_2, n371_2, n372_2, n373_2, n374_2, \inst_line_buf/r_mipi_rx_data_1P[0]_2 , 
        \inst_line_buf/r_mipi_rx_valid_1P_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 , 
        \inst_line_buf/r_mipi_rx_hsync_2P , \inst_line_buf/r_mipi_tx_x_1P[0]_2 , 
        \inst_line_buf/r_mipi_rx_full_1P_2 , \inst_line_buf/r_mipi_tx_en_1P , 
        \inst_line_buf/r_mipi_tx_x_inc_1P , \inst_line_buf/r_mipi_tx_b_1P[0] , 
        \inst_line_buf/r_mipi_tx_data_4P[0] , \inst_line_buf/r_mipi_tx_hsync_1P_2 , 
        \inst_line_buf/r_mipi_tx_valid_1P_2 , \inst_line_buf/r_mipi_tx_hsync_2P_2 , 
        \inst_line_buf/r_mipi_tx_valid_2P_2 , \inst_line_buf/r_mipi_tx_hsync_3P_2 , 
        \inst_line_buf/r_mipi_tx_valid_3P_2 , \inst_line_buf/r_mipi_tx_hsync_4P_2 , 
        \inst_line_buf/r_mipi_tx_valid_4P_2 , n394, n395, \inst_line_buf/r_mipi_tx_hsync_5P_2 , 
        \inst_line_buf/r_mipi_tx_valid_5P_2 , \inst_line_buf/r_mipi_rx_hsync_1P , 
        n401, n402, n403, n404, n405, n406, n407, n408, n409, 
        n410, n411, n412, n413, n414, n415, n416, n417, n418, 
        n419, n420, n421, n422, n423, n424, \inst_line_buf/r_mipi_rx_data_1P[1]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[2]_2 , \inst_line_buf/r_mipi_rx_data_1P[3]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[4]_2 , \inst_line_buf/r_mipi_rx_data_1P[5]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[6]_2 , \inst_line_buf/r_mipi_rx_data_1P[7]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[8]_2 , \inst_line_buf/r_mipi_rx_data_1P[9]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[10]_2 , \inst_line_buf/r_mipi_rx_data_1P[11]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[12]_2 , \inst_line_buf/r_mipi_rx_data_1P[13]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[14]_2 , \inst_line_buf/r_mipi_rx_data_1P[15]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[16]_2 , \inst_line_buf/r_mipi_rx_data_1P[17]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[18]_2 , \inst_line_buf/r_mipi_rx_data_1P[19]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[20]_2 , \inst_line_buf/r_mipi_rx_data_1P[21]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[22]_2 , \inst_line_buf/r_mipi_rx_data_1P[23]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[24]_2 , \inst_line_buf/r_mipi_rx_data_1P[25]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[26]_2 , \inst_line_buf/r_mipi_rx_data_1P[27]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[28]_2 , \inst_line_buf/r_mipi_rx_data_1P[29]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[30]_2 , \inst_line_buf/r_mipi_rx_data_1P[31]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[32]_2 , \inst_line_buf/r_mipi_rx_data_1P[33]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[34]_2 , \inst_line_buf/r_mipi_rx_data_1P[35]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[36]_2 , \inst_line_buf/r_mipi_rx_data_1P[37]_2 , 
        \inst_line_buf/r_mipi_rx_data_1P[38]_2 , \inst_line_buf/r_mipi_rx_data_1P[39]_2 , 
        \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
        \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
        \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
        \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
        \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
        \inst_line_buf/r_mipi_tx_x_1P[1]_2 , \inst_line_buf/r_mipi_tx_x_1P[2]_2 , 
        \inst_line_buf/r_mipi_tx_x_1P[3]_2 , \inst_line_buf/r_mipi_tx_x_1P[4]_2 , 
        \inst_line_buf/r_mipi_tx_x_1P[5]_2 , \inst_line_buf/r_mipi_tx_x_1P[6]_2 , 
        \inst_line_buf/r_mipi_tx_x_1P[7]_2 , \inst_line_buf/r_mipi_tx_x_1P[8]_2 , 
        \inst_line_buf/r_mipi_tx_x_1P[9]_2 , \inst_line_buf/r_mipi_tx_x_1P[10]_2 , 
        \inst_line_buf/r_mipi_tx_b_1P[1] , \inst_line_buf/r_mipi_tx_b_1P[2] , 
        \inst_line_buf/r_mipi_tx_data_4P[1] , \inst_line_buf/r_mipi_tx_data_4P[2] , 
        \inst_line_buf/r_mipi_tx_data_4P[3] , \inst_line_buf/r_mipi_tx_data_4P[4] , 
        \inst_line_buf/r_mipi_tx_data_4P[5] , \inst_line_buf/r_mipi_tx_data_4P[6] , 
        \inst_line_buf/r_mipi_tx_data_4P[7] , \inst_line_buf/r_mipi_tx_data_4P[8] , 
        \inst_line_buf/r_mipi_tx_data_4P[9] , \inst_line_buf/r_mipi_tx_data_4P[10] , 
        \inst_line_buf/r_mipi_tx_data_4P[11] , \inst_line_buf/r_mipi_tx_data_4P[12] , 
        \inst_line_buf/r_mipi_tx_data_4P[13] , \inst_line_buf/r_mipi_tx_data_4P[14] , 
        \inst_line_buf/r_mipi_tx_data_4P[15] , \inst_line_buf/r_mipi_tx_data_4P[16] , 
        \inst_line_buf/r_mipi_tx_data_4P[17] , \inst_line_buf/r_mipi_tx_data_4P[18] , 
        \inst_line_buf/r_mipi_tx_data_4P[19] , \inst_line_buf/r_mipi_tx_data_4P[20] , 
        \inst_line_buf/r_mipi_tx_data_4P[21] , \inst_line_buf/r_mipi_tx_data_4P[22] , 
        \inst_line_buf/r_mipi_tx_data_4P[23] , \inst_line_buf/r_mipi_tx_data_4P[24] , 
        \inst_line_buf/r_mipi_tx_data_4P[25] , \inst_line_buf/r_mipi_tx_data_4P[26] , 
        \inst_line_buf/r_mipi_tx_data_4P[27] , \inst_line_buf/r_mipi_tx_data_4P[28] , 
        \inst_line_buf/r_mipi_tx_data_4P[29] , \inst_line_buf/r_mipi_tx_data_4P[30] , 
        \inst_line_buf/r_mipi_tx_data_4P[31] , \inst_line_buf/r_mipi_tx_data_4P[32] , 
        \inst_line_buf/r_mipi_tx_data_4P[33] , \inst_line_buf/r_mipi_tx_data_4P[34] , 
        \inst_line_buf/r_mipi_tx_data_4P[35] , \inst_line_buf/r_mipi_tx_data_4P[36] , 
        \inst_line_buf/r_mipi_tx_data_4P[37] , \inst_line_buf/r_mipi_tx_data_4P[38] , 
        \inst_line_buf/r_mipi_tx_data_4P[39] , \inst_line_buf/r_mipi_tx_data_4P[40] , 
        \inst_line_buf/r_mipi_tx_data_4P[41] , \inst_line_buf/r_mipi_tx_data_4P[42] , 
        \inst_line_buf/r_mipi_tx_data_4P[43] , \inst_line_buf/r_mipi_tx_data_4P[44] , 
        \inst_line_buf/r_mipi_tx_data_4P[45] , \inst_line_buf/r_mipi_tx_data_4P[46] , 
        \inst_line_buf/r_mipi_tx_data_4P[47] , \inst_line_buf/r_mipi_tx_data_4P[48] , 
        \inst_line_buf/r_mipi_tx_data_4P[49] , \inst_line_buf/r_mipi_tx_data_4P[50] , 
        \inst_line_buf/r_mipi_tx_data_4P[51] , \inst_line_buf/r_mipi_tx_data_4P[52] , 
        \inst_line_buf/r_mipi_tx_data_4P[53] , \inst_line_buf/r_mipi_tx_data_4P[54] , 
        \inst_line_buf/r_mipi_tx_data_4P[55] , \inst_line_buf/r_mipi_tx_data_4P[56] , 
        \inst_line_buf/r_mipi_tx_data_4P[57] , \inst_line_buf/r_mipi_tx_data_4P[58] , 
        \inst_line_buf/r_mipi_tx_data_4P[59] , \inst_line_buf/r_mipi_tx_data_4P[60] , 
        \inst_line_buf/r_mipi_tx_data_4P[61] , \inst_line_buf/r_mipi_tx_data_4P[62] , 
        \inst_line_buf/r_mipi_tx_data_4P[63] , \inst_line_buf/r_mipi_tx_data_4P[64] , 
        \inst_line_buf/r_mipi_tx_data_4P[65] , \inst_line_buf/r_mipi_tx_data_4P[66] , 
        \inst_line_buf/r_mipi_tx_data_4P[67] , \inst_line_buf/r_mipi_tx_data_4P[68] , 
        \inst_line_buf/r_mipi_tx_data_4P[69] , \inst_line_buf/r_mipi_tx_data_4P[70] , 
        \inst_line_buf/r_mipi_tx_data_4P[71] , \inst_line_buf/r_mipi_tx_data_4P[72] , 
        \inst_line_buf/r_mipi_tx_data_4P[73] , \inst_line_buf/r_mipi_tx_data_4P[74] , 
        \inst_line_buf/r_mipi_tx_data_4P[75] , \inst_line_buf/r_mipi_tx_data_4P[76] , 
        \inst_line_buf/r_mipi_tx_data_4P[77] , \inst_line_buf/r_mipi_tx_data_4P[78] , 
        \inst_line_buf/r_mipi_tx_data_4P[79] , \inst_line_buf/r_mipi_tx_data_4P[80] , 
        \inst_line_buf/r_mipi_tx_data_4P[81] , \inst_line_buf/r_mipi_tx_data_4P[82] , 
        \inst_line_buf/r_mipi_tx_data_4P[83] , \inst_line_buf/r_mipi_tx_data_4P[84] , 
        \inst_line_buf/r_mipi_tx_data_4P[85] , \inst_line_buf/r_mipi_tx_data_4P[86] , 
        \inst_line_buf/r_mipi_tx_data_4P[87] , \inst_line_buf/r_mipi_tx_data_4P[88] , 
        \inst_line_buf/r_mipi_tx_data_4P[89] , \inst_line_buf/r_mipi_tx_data_4P[90] , 
        \inst_line_buf/r_mipi_tx_data_4P[91] , \inst_line_buf/r_mipi_tx_data_4P[92] , 
        \inst_line_buf/r_mipi_tx_data_4P[93] , \inst_line_buf/r_mipi_tx_data_4P[94] , 
        \inst_line_buf/r_mipi_tx_data_4P[95] , \inst_line_buf/r_mipi_tx_data_4P[96] , 
        \inst_line_buf/r_mipi_tx_data_4P[97] , \inst_line_buf/r_mipi_tx_data_4P[98] , 
        \inst_line_buf/r_mipi_tx_data_4P[99] , \inst_line_buf/r_mipi_tx_data_4P[100] , 
        \inst_line_buf/r_mipi_tx_data_4P[101] , \inst_line_buf/r_mipi_tx_data_4P[102] , 
        \inst_line_buf/r_mipi_tx_data_4P[103] , \inst_line_buf/r_mipi_tx_data_4P[104] , 
        \inst_line_buf/r_mipi_tx_data_4P[105] , \inst_line_buf/r_mipi_tx_data_4P[106] , 
        \inst_line_buf/r_mipi_tx_data_4P[107] , \inst_line_buf/r_mipi_tx_data_4P[108] , 
        \inst_line_buf/r_mipi_tx_data_4P[109] , \inst_line_buf/r_mipi_tx_data_4P[110] , 
        \inst_line_buf/r_mipi_tx_data_4P[111] , \inst_line_buf/r_mipi_tx_data_4P[112] , 
        \inst_line_buf/r_mipi_tx_data_4P[113] , \inst_line_buf/r_mipi_tx_data_4P[114] , 
        \inst_line_buf/r_mipi_tx_data_4P[115] , \inst_line_buf/r_mipi_tx_data_4P[116] , 
        \inst_line_buf/r_mipi_tx_data_4P[117] , \inst_line_buf/r_mipi_tx_data_4P[118] , 
        \inst_line_buf/r_mipi_tx_data_4P[119] , \inst_line_buf/r_mipi_tx_data_5P[60] , 
        \inst_line_buf/r_mipi_tx_data_5P[61] , \inst_line_buf/r_mipi_tx_data_5P[62] , 
        \inst_line_buf/r_mipi_tx_data_5P[63] , \inst_line_buf/r_mipi_tx_data_5P[64] , 
        \inst_line_buf/r_mipi_tx_data_5P[65] , \inst_line_buf/r_mipi_tx_data_5P[66] , 
        \inst_line_buf/r_mipi_tx_data_5P[67] , \inst_line_buf/r_mipi_tx_data_5P[68] , 
        \inst_line_buf/r_mipi_tx_data_5P[69] , \inst_line_buf/r_mipi_tx_data_5P[70] , 
        \inst_line_buf/r_mipi_tx_data_5P[71] , \inst_line_buf/r_mipi_tx_data_5P[72] , 
        \inst_line_buf/r_mipi_tx_data_5P[73] , \inst_line_buf/r_mipi_tx_data_5P[74] , 
        \inst_line_buf/r_mipi_tx_data_5P[75] , \inst_line_buf/r_mipi_tx_data_5P[76] , 
        \inst_line_buf/r_mipi_tx_data_5P[77] , \inst_line_buf/r_mipi_tx_data_5P[78] , 
        \inst_line_buf/r_mipi_tx_data_5P[79] , \inst_line_buf/r_mipi_tx_data_5P[80] , 
        \inst_line_buf/r_mipi_tx_data_5P[81] , \inst_line_buf/r_mipi_tx_data_5P[82] , 
        \inst_line_buf/r_mipi_tx_data_5P[83] , \inst_line_buf/r_mipi_tx_data_5P[84] , 
        \inst_line_buf/r_mipi_tx_data_5P[85] , \inst_line_buf/r_mipi_tx_data_5P[86] , 
        \inst_line_buf/r_mipi_tx_data_5P[87] , \inst_line_buf/r_mipi_tx_data_5P[88] , 
        \inst_line_buf/r_mipi_tx_data_5P[89] , \inst_line_buf/r_mipi_tx_data_5P[90] , 
        \inst_line_buf/r_mipi_tx_data_5P[91] , \inst_line_buf/r_mipi_tx_data_5P[92] , 
        \inst_line_buf/r_mipi_tx_data_5P[93] , \inst_line_buf/r_mipi_tx_data_5P[94] , 
        \inst_line_buf/r_mipi_tx_data_5P[95] , \inst_line_buf/r_mipi_tx_data_5P[96] , 
        \inst_line_buf/r_mipi_tx_data_5P[97] , \inst_line_buf/r_mipi_tx_data_5P[98] , 
        \inst_line_buf/r_mipi_tx_data_5P[99] , \inst_line_buf/r_mipi_tx_data_5P[100] , 
        \inst_line_buf/r_mipi_tx_data_5P[101] , \inst_line_buf/r_mipi_tx_data_5P[102] , 
        \inst_line_buf/r_mipi_tx_data_5P[103] , \inst_line_buf/r_mipi_tx_data_5P[104] , 
        \inst_line_buf/r_mipi_tx_data_5P[105] , \inst_line_buf/r_mipi_tx_data_5P[106] , 
        \inst_line_buf/r_mipi_tx_data_5P[107] , \inst_line_buf/r_mipi_tx_data_5P[108] , 
        \inst_line_buf/r_mipi_tx_data_5P[109] , \inst_line_buf/r_mipi_tx_data_5P[110] , 
        \inst_line_buf/r_mipi_tx_data_5P[111] , \inst_line_buf/r_mipi_tx_data_5P[112] , 
        \inst_line_buf/r_mipi_tx_data_5P[113] , \inst_line_buf/r_mipi_tx_data_5P[114] , 
        \inst_line_buf/r_mipi_tx_data_5P[115] , \inst_line_buf/r_mipi_tx_data_5P[116] , 
        \inst_line_buf/r_mipi_tx_data_5P[117] , \inst_line_buf/r_mipi_tx_data_5P[118] , 
        \inst_line_buf/r_mipi_tx_data_5P[119] , \inst_line_buf/w_mipi_tx_data_3P[0] , 
        \inst_dly/n28 , \inst_line_buf/w_mipi_tx_data_3P[1] , \inst_line_buf/w_mipi_tx_data_3P[2] , 
        \inst_line_buf/w_mipi_tx_data_3P[3] , \inst_line_buf/w_mipi_tx_data_3P[4] , 
        \inst_line_buf/w_mipi_tx_data_3P[5] , \inst_line_buf/w_mipi_tx_data_3P[6] , 
        \inst_line_buf/w_mipi_tx_data_3P[7] , \inst_line_buf/w_mipi_tx_data_3P[8] , 
        \inst_line_buf/w_mipi_tx_data_3P[9] , \inst_line_buf/w_mipi_tx_data_3P[10] , 
        \inst_line_buf/w_mipi_tx_data_3P[11] , \inst_line_buf/w_mipi_tx_data_3P[12] , 
        \inst_line_buf/w_mipi_tx_data_3P[13] , \inst_line_buf/w_mipi_tx_data_3P[14] , 
        \inst_line_buf/w_mipi_tx_data_3P[15] , \inst_line_buf/w_mipi_tx_data_3P[16] , 
        \inst_line_buf/w_mipi_tx_data_3P[17] , \inst_line_buf/w_mipi_tx_data_3P[18] , 
        \inst_line_buf/w_mipi_tx_data_3P[19] , \inst_line_buf/w_mipi_tx_data_3P[20] , 
        \inst_line_buf/w_mipi_tx_data_3P[21] , \inst_line_buf/w_mipi_tx_data_3P[22] , 
        \inst_line_buf/w_mipi_tx_data_3P[23] , \inst_line_buf/w_mipi_tx_data_3P[24] , 
        \inst_line_buf/w_mipi_tx_data_3P[25] , \inst_line_buf/w_mipi_tx_data_3P[26] , 
        \inst_line_buf/w_mipi_tx_data_3P[27] , \inst_line_buf/w_mipi_tx_data_3P[28] , 
        \inst_line_buf/w_mipi_tx_data_3P[29] , \inst_line_buf/w_mipi_tx_data_3P[30] , 
        \inst_line_buf/w_mipi_tx_data_3P[31] , \inst_line_buf/w_mipi_tx_data_3P[32] , 
        \inst_line_buf/w_mipi_tx_data_3P[33] , \inst_line_buf/w_mipi_tx_data_3P[34] , 
        \inst_line_buf/w_mipi_tx_data_3P[35] , \inst_line_buf/w_mipi_tx_data_3P[36] , 
        \inst_line_buf/w_mipi_tx_data_3P[37] , \inst_line_buf/w_mipi_tx_data_3P[38] , 
        \inst_line_buf/w_mipi_tx_data_3P[39] , \mipi_pclk~O , n2442, n2441, 
        n2440, n2439, n2438, n2437, n2436, n2435, n2434, n2433, 
        n2432, n2431, n2430, n2429, n2428, n2427, n2426, n2425, 
        n805, n806, n807, n808, n809, n810, n811, n812, n813, 
        n814, n815, n816, n817, n818, n819, n820, n821, n822, 
        n823, n824, n825, n826, n827, n828, n829, n830, n831, 
        n832, n833, n834, n835, n836, n837, n838, n839, n840, 
        n841, n842, n843, n844, n845, n846, n847, n848, n849, 
        n850, n851, n852, n853, n854, n855, n856, n857, n858, 
        n859, n860, n861, n862, n863, n864, n865, n866, n867, 
        n868, n869, n870, n871, n872, n873, n874_2, n875_2, 
        n876, n877, n878, n879, n880, n881, n882, n883, n884, 
        n885_2, n886, n887, n888, n889, n890_2, n891, n892, 
        n893, n894, n895_2, n896, n897, n898, n899, n900_2, 
        n901, n902, n903, n904, n905_2, n906, n907, n908, n909, 
        n910_2, n911, n912, n913, n914, n915_2, n916, n917, 
        n918, n919, n920_2, n921, n922, n923, n924, n925_2, 
        n926, n927, n928, n929, n930_2, n931, n932, n933, n934, 
        n935_2, n936, n937, n938, n939, n940_2, n941, n942, 
        n943, n944, n945_2, n946, n947, n948, n949, n950_2, 
        n951, n952, n953, n954, n955_2, n956, n957, n958, n959, 
        n960, n961, n962, n963, n964, n965, n966, n967, n968, 
        n969, n970, n971, n972, n973, n974, n975, n976, n977, 
        n978, n979, n980, \r_raddr_1P[1]_2 , \r_raddr_1P[2]_2 , \r_raddr_1P[3]_2 , 
        \r_raddr_1P[4]_2 , \r_raddr_1P[5]_2 , \r_raddr_1P[6]_2 , \r_raddr_1P[7]_2 , 
        \r_raddr_1P[8]_2 , \r_raddr_1P[9]_2 , \r_raddr_1P[10]_2 , \r_raddr_1P[11]_2 , 
        \r_raddr_1P[12]_2 , \inst_dly/n29 , n995, n996, \inst_dly/n24 , 
        n998, n999, n1000, n1001, n1026, n1027, n1028, n1029, 
        n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, 
        n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
        n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
        n1054, n1055, n1056, n1057, n1058, n1059, n1060_2, n1061, 
        n1062, n1063, n1065_2, n1066, n1067, n1068, n1071, n1072, 
        n1073, n1074, n1075_2, n1076, n1077, n1078, n1079, n1080_2, 
        n1081, n1082, n1083, n1084, n1085_2, n1086, n1087, n1088, 
        n1089, n1090_2, n1091, n271, n874, n1247, n1251, n1254, 
        n1261, n380, ceg_net83, \equal_59/n31 , n875, n1272, n1277, 
        n1280, n1282, n1288, n885, n890, n895, n900, n905, n910, 
        n915, n920, n925, n930, n935, n940, n945, n950, n955, 
        n1309, n1312, n1315, n1318, n379, n378, n377, n376, 
        n375, n374, n373, n372, n371, n370, n369, n368, n367, 
        n366, n365, n390, n389, n1482, n1484, n1490, n1498, 
        n1501, n1506, \inst_line_buf/even_line_pix_0[0] , \inst_line_buf/n1296 , 
        ceg_net98, \inst_line_buf/n1381 , ceg_net101, \inst_line_buf/n2531 , 
        ceg_net104, \inst_line_buf/n1385 , ceg_net140, \inst_line_buf/n1387 , 
        \inst_line_buf/n1510 , n1533, n1548, n1550, n1553, n1555, 
        \inst_line_buf/odd_line_pix_0[1] , \inst_line_buf/odd_line_pix_0[2] , 
        \inst_line_buf/odd_line_pix_0[3] , \inst_line_buf/odd_line_pix_0[4] , 
        \inst_line_buf/odd_line_pix_0[5] , \inst_line_buf/odd_line_pix_0[6] , 
        \inst_line_buf/odd_line_pix_0[7] , \inst_line_buf/odd_line_pix_0[8] , 
        \inst_line_buf/odd_line_pix_0[9] , \inst_line_buf/mipi_inst1_DATA_filtered[10] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[11] , \inst_line_buf/mipi_inst1_DATA_filtered[12] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[13] , \inst_line_buf/mipi_inst1_DATA_filtered[14] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[15] , \inst_line_buf/mipi_inst1_DATA_filtered[16] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[17] , \inst_line_buf/mipi_inst1_DATA_filtered[18] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[19] , \inst_line_buf/even_line_pix_2[0] , 
        \inst_line_buf/odd_line_pix_2[1] , \inst_line_buf/odd_line_pix_2[2] , 
        \inst_line_buf/odd_line_pix_2[3] , \inst_line_buf/odd_line_pix_2[4] , 
        \inst_line_buf/odd_line_pix_2[5] , \inst_line_buf/odd_line_pix_2[6] , 
        \inst_line_buf/odd_line_pix_2[7] , \inst_line_buf/odd_line_pix_2[8] , 
        \inst_line_buf/odd_line_pix_2[9] , \inst_line_buf/mipi_inst1_DATA_filtered[30] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[31] , \inst_line_buf/mipi_inst1_DATA_filtered[32] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[33] , \inst_line_buf/mipi_inst1_DATA_filtered[34] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[35] , \inst_line_buf/mipi_inst1_DATA_filtered[36] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[37] , \inst_line_buf/mipi_inst1_DATA_filtered[38] , 
        \inst_line_buf/mipi_inst1_DATA_filtered[39] , \inst_line_buf/n1295 , 
        \inst_line_buf/n1294 , \inst_line_buf/n1293 , \inst_line_buf/n1292 , 
        \inst_line_buf/n1291 , \inst_line_buf/n1290 , \inst_line_buf/n1289 , 
        \inst_line_buf/n1288 , \inst_line_buf/n1287 , \inst_line_buf/n1283 , 
        \inst_line_buf/n1380 , \inst_line_buf/n1379 , \inst_line_buf/n1378 , 
        \inst_line_buf/n1377 , \inst_line_buf/n1376 , \inst_line_buf/n1375 , 
        \inst_line_buf/n1374 , \inst_line_buf/n1373 , \inst_line_buf/n1372 , 
        \inst_line_buf/n1384 , \inst_line_buf/n1383 , \inst_line_buf/n1509 , 
        \inst_line_buf/n1508 , \inst_line_buf/n1507 , \inst_line_buf/n1506 , 
        \inst_line_buf/n1505 , \inst_line_buf/n1504 , \inst_line_buf/n1503 , 
        \inst_line_buf/n1502 , \inst_line_buf/n1501 , \inst_line_buf/n1500 , 
        \inst_line_buf/n1499 , \inst_line_buf/n1498 , \inst_line_buf/n1497 , 
        \inst_line_buf/n1496 , \inst_line_buf/n1495 , \inst_line_buf/n1494 , 
        \inst_line_buf/n1493 , \inst_line_buf/n1492 , \inst_line_buf/n1491 , 
        \inst_line_buf/n1490 , \inst_line_buf/n1489 , \inst_line_buf/n1488 , 
        \inst_line_buf/n1487 , \inst_line_buf/n1486 , \inst_line_buf/n1485 , 
        \inst_line_buf/n1484 , \inst_line_buf/n1483 , \inst_line_buf/n1482 , 
        \inst_line_buf/n1481 , \inst_line_buf/n1480 , \inst_line_buf/n1479 , 
        \inst_line_buf/n1478 , \inst_line_buf/n1477 , \inst_line_buf/n1476 , 
        \inst_line_buf/n1475 , \inst_line_buf/n1474 , \inst_line_buf/n1473 , 
        \inst_line_buf/n1472 , \inst_line_buf/n1471 , \inst_line_buf/n1470 , 
        \inst_line_buf/n1469 , \inst_line_buf/n1468 , \inst_line_buf/n1467 , 
        \inst_line_buf/n1466 , \inst_line_buf/n1465 , \inst_line_buf/n1464 , 
        \inst_line_buf/n1463 , \inst_line_buf/n1462 , \inst_line_buf/n1461 , 
        \inst_line_buf/n1460 , \inst_line_buf/n1459 , \inst_line_buf/n1458 , 
        \inst_line_buf/n1457 , \inst_line_buf/n1456 , \inst_line_buf/n1455 , 
        \inst_line_buf/n1454 , \inst_line_buf/n1453 , \inst_line_buf/n1452 , 
        \inst_line_buf/n1451 , \inst_line_buf/n1450 , \inst_line_buf/n1449 , 
        \inst_line_buf/n1448 , \inst_line_buf/n1447 , \inst_line_buf/n1446 , 
        \inst_line_buf/n1445 , \inst_line_buf/n1444 , \inst_line_buf/n1443 , 
        \inst_line_buf/n1442 , \inst_line_buf/n1441 , \inst_line_buf/n1440 , 
        \inst_line_buf/n1439 , \inst_line_buf/n1438 , \inst_line_buf/n1437 , 
        \inst_line_buf/n1436 , \inst_line_buf/n1435 , \inst_line_buf/n1434 , 
        \inst_line_buf/n1433 , \inst_line_buf/n1432 , \inst_line_buf/n1431 , 
        \inst_line_buf/n1430 , \inst_line_buf/n1429 , \inst_line_buf/n1428 , 
        \inst_line_buf/n1427 , \inst_line_buf/n1426 , \inst_line_buf/n1425 , 
        \inst_line_buf/n1424 , \inst_line_buf/n1423 , \inst_line_buf/n1422 , 
        \inst_line_buf/n1421 , \inst_line_buf/n1420 , \inst_line_buf/n1419 , 
        \inst_line_buf/n1418 , \inst_line_buf/n1417 , \inst_line_buf/n1416 , 
        \inst_line_buf/n1415 , \inst_line_buf/n1414 , \inst_line_buf/n1413 , 
        \inst_line_buf/n1412 , \inst_line_buf/n1411 , \inst_line_buf/n1410 , 
        \inst_line_buf/n1409 , \inst_line_buf/n1408 , \inst_line_buf/n1407 , 
        \inst_line_buf/n1406 , \inst_line_buf/n1405 , \inst_line_buf/n1404 , 
        \inst_line_buf/n1403 , \inst_line_buf/n1402 , \inst_line_buf/n1401 , 
        \inst_line_buf/n1400 , \inst_line_buf/n1399 , \inst_line_buf/n1398 , 
        \inst_line_buf/n1397 , \inst_line_buf/n1396 , \inst_line_buf/n1395 , 
        \inst_line_buf/n1394 , \inst_line_buf/n1393 , \inst_line_buf/n1392 , 
        \inst_line_buf/n1391 , n1502, n2071, n2074, n2077, n2080, 
        n2083, n2086, n2089, n2092, n2094, n2096, n2098, n2100, 
        n2102, n2104, n2106, n2115, n2118, n2121, n2124, n2127, 
        n2130, n2133, n2136, n2139, n2142, n2146, n2148, n2150, 
        n2152, n2154, n2156, n2159, n2161, n2163, n2165, n2167, 
        n2169, n2171, n2173, n1060, n1065, n1070, n1075, n1080, 
        n1085, n1090, n1095, n1100, n1105, n1110, n1115, n1504, 
        \inst_dly/r_rdata_1P[0] , n2221, n2223, n2278, n2281, n2284, 
        n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, 
        n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, 
        n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, 
        n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, 
        n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, 
        n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
        n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, 
        n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, 
        n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, 
        n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, 
        n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, 
        n2418, n2419, n2420, n2421, n2422, n2423, n2424;
    
    assign mipi_inst1_DPHY_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_VC_ENA[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_VC_ENA[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_VC_ENA[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_VC_ENA[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_LANES[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_LANES[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst1_CLEAR = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign standby = mipi_inst1_HSYNC[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign rx_status = mipi_inst1_VSYNC[0] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign rx_status2 = mipi_inst1_ERR[9] /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_INPUT=TRUE */ ;
    assign mipi_inst2_DPHY_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_RSTN = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HSYNC = rx_status3 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_DATA[63] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_DATA[62] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_DATA[61] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_DATA[60] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_TYPE[5] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_TYPE[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_TYPE[3] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_TYPE[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_TYPE[1] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_TYPE[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_LANES[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_LANES[0] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_FRAME_MODE = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[15] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[14] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[13] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[12] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[11] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[10] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[9] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[8] = 1'b1 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[6] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[5] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[4] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_VC[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_VC[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_ENTER[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_ENTER[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_ENTER[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_ENTER[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_EXIT[3] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_EXIT[2] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_EXIT[1] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_EXIT[0] = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_CLK_ENTER = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_ULPS_CLK_EXIT = 1'b0 /* verific EFX_ATTRIBUTE_PORT__IS_PRIMARY_OUTPUT=TRUE */ ;
    assign mipi_inst2_HRES[7] = 1'b1 /* verific EFX_ATTRIBUTE_CELL_NAME=VCC */ ;
    assign mipi_inst2_HRES[2] = 1'b0 /* verific EFX_ATTRIBUTE_CELL_NAME=GND */ ;
    EFX_LUT4 LUT__3516 (.I0(n2330), .I1(\key1_counter[4] ), .I2(\key1_counter[5] ), 
            .I3(\key1_counter[6] ), .O(n2331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__3516.LUTMASK = 16'hf400;
    EFX_FF \r_mipi_rx_data_1P[35]~FF  (.D(mipi_inst1_DATA[35]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[35]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[35]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[35]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[35]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[35]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[35]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[34]~FF  (.D(mipi_inst1_DATA[34]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[34]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[34]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[34]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[34]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[34]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[34]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[21]~FF  (.D(mipi_inst1_DATA[21]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[21]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[21]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[21]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[21]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[21]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[21]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[20]~FF  (.D(mipi_inst1_DATA[20]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[20]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[20]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[20]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[20]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[20]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[20]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[39]~FF  (.D(mipi_inst1_DATA[39]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[39]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[39]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[39]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[39]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[39]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[39]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[38]~FF  (.D(mipi_inst1_DATA[38]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[38]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[38]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[38]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[38]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[38]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[38]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[37]~FF  (.D(mipi_inst1_DATA[37]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[37]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[37]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[37]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[37]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[37]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[37]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[36]~FF  (.D(mipi_inst1_DATA[36]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[36]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[36]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[36]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[36]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[36]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[36]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[19]~FF  (.D(mipi_inst1_DATA[19]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[19]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[19]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[19]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[19]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[19]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[19]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[18]~FF  (.D(mipi_inst1_DATA[18]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[18]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[18]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[18]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[18]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[18]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[18]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[17]~FF  (.D(mipi_inst1_DATA[17]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[17]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[17]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[17]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[17]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[17]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[17]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[16]~FF  (.D(mipi_inst1_DATA[16]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[16]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[16]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[16]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[16]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[16]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[16]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[15]~FF  (.D(mipi_inst1_DATA[15]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[15]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[15]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[15]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[15]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[15]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[15]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[14]~FF  (.D(mipi_inst1_DATA[14]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[14]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[14]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[14]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[14]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[14]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[14]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[13]~FF  (.D(mipi_inst1_DATA[13]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[13]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[13]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[13]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[13]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[13]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[13]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[12]~FF  (.D(mipi_inst1_DATA[12]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[12]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[12]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[12]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[12]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[12]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[11]~FF  (.D(mipi_inst1_DATA[11]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[11]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[11]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[11]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[11]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[11]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[23]~FF  (.D(mipi_inst1_DATA[23]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[23]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[23]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[23]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[23]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[23]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[23]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[10]~FF  (.D(mipi_inst1_DATA[10]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[10]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[10]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[10]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[10]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[10]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[9]~FF  (.D(mipi_inst1_DATA[9]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[9]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[8]~FF  (.D(mipi_inst1_DATA[8]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[8]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[7]~FF  (.D(mipi_inst1_DATA[7]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[22]~FF  (.D(mipi_inst1_DATA[22]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[22]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[22]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[22]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[22]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[22]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[22]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[6]~FF  (.D(mipi_inst1_DATA[6]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[5]~FF  (.D(mipi_inst1_DATA[5]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[4]~FF  (.D(mipi_inst1_DATA[4]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[4]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[3]~FF  (.D(mipi_inst1_DATA[3]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[3]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[2]~FF  (.D(mipi_inst1_DATA[2]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[2]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[1]~FF  (.D(mipi_inst1_DATA[1]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[1]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[33]~FF  (.D(mipi_inst1_DATA[33]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[33]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[33]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[33]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[33]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[33]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[33]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[0]~FF  (.D(mipi_inst1_DATA[0]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[0]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[32]~FF  (.D(mipi_inst1_DATA[32]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[32]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[32]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[32]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[32]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[32]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[32]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[31]~FF  (.D(mipi_inst1_DATA[31]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[31]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[31]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[31]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[31]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[31]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[31]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_valid_1P~FF  (.D(mipi_inst1_VALID), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(r_mipi_rx_valid_1P_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_valid_1P~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_valid_1P~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_valid_1P~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_valid_1P~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_valid_1P~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_valid_1P~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_valid_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[0]_2~FF  (.D(\key1_counter[0]_2 ), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[0]_2~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[0]_2~FF .D_POLARITY = 1'b0;
    defparam \key1_counter[0]_2~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[0]_2~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[30]~FF  (.D(mipi_inst1_DATA[30]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[30]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[30]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[30]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[30]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[30]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[30]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[29]~FF  (.D(mipi_inst1_DATA[29]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[29]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[29]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[29]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[29]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[29]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[29]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[28]~FF  (.D(mipi_inst1_DATA[28]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[28]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[28]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[28]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[28]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[28]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[28]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[0]~FF  (.D(n380), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[0]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[0]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[0]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[0]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[0]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[0]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[25]~FF  (.D(mipi_inst1_DATA[25]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[25]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[25]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[25]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[25]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[25]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[25]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[24]~FF  (.D(mipi_inst1_DATA[24]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[24]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[24]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[24]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[24]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[24]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[24]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \red_gain[0]~FF  (.D(\red_gain[0] ), .CE(\equal_59/n31 ), .CLK(\mipi_pclk~O ), 
           .SR(n875), .Q(\red_gain[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \red_gain[0]~FF .CLK_POLARITY = 1'b1;
    defparam \red_gain[0]~FF .CE_POLARITY = 1'b0;
    defparam \red_gain[0]~FF .SR_POLARITY = 1'b1;
    defparam \red_gain[0]~FF .D_POLARITY = 1'b0;
    defparam \red_gain[0]~FF .SR_SYNC = 1'b1;
    defparam \red_gain[0]~FF .SR_VALUE = 1'b0;
    defparam \red_gain[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[0]_2~FF  (.D(\r_waddr_1P[0]_2 ), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[0]_2~FF .D_POLARITY = 1'b0;
    defparam \r_waddr_1P[0]_2~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[0]_2~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[27]~FF  (.D(mipi_inst1_DATA[27]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[27]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[27]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[27]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[27]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[27]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[27]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_data_1P[26]~FF  (.D(mipi_inst1_DATA[26]), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_mipi_rx_data_1P[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_data_1P[26]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[26]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[26]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_data_1P[26]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_data_1P[26]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_data_1P[26]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_data_1P[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[0]_2~FF  (.D(\r_raddr_1P[0]_2 ), .CE(r_rden_1P_2), 
           .CLK(\mipi_pclk~O ), .SR(i_arstn), .Q(\r_raddr_1P[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[0]_2~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[0]_2~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[0]_2~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[0]_2~FF .D_POLARITY = 1'b0;
    defparam \r_raddr_1P[0]_2~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[0]_2~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[0]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_rden_1P~FF  (.D(1'b1), .CE(\r_waddr_1P[10]_2 ), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(r_rden_1P_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_rden_1P~FF .CLK_POLARITY = 1'b1;
    defparam \r_rden_1P~FF .CE_POLARITY = 1'b1;
    defparam \r_rden_1P~FF .SR_POLARITY = 1'b0;
    defparam \r_rden_1P~FF .D_POLARITY = 1'b1;
    defparam \r_rden_1P~FF .SR_SYNC = 1'b0;
    defparam \r_rden_1P~FF .SR_VALUE = 1'b0;
    defparam \r_rden_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_mipi_rx_hsync_1P[0]~FF  (.D(standby), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_mipi_rx_hsync_1P[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(157)
    defparam \r_mipi_rx_hsync_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \r_mipi_rx_hsync_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \r_mipi_rx_hsync_1P[0]~FF .SR_POLARITY = 1'b0;
    defparam \r_mipi_rx_hsync_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \r_mipi_rx_hsync_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \r_mipi_rx_hsync_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \r_mipi_rx_hsync_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[1]~FF  (.D(n885), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[1]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[2]~FF  (.D(n890), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[2]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[3]~FF  (.D(n895), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[3]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[4]~FF  (.D(n900), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[4]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[5]~FF  (.D(n905), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[5]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[6]~FF  (.D(n910), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[6]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[7]~FF  (.D(n915), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[7]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[8]~FF  (.D(n920), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[8]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[9]~FF  (.D(n925), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[9]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[10]~FF  (.D(n930), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[10]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[10]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[11]~FF  (.D(n935), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[11]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[11]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[12]~FF  (.D(n940), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[12]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[12]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[13]~FF  (.D(n945), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[13]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[13]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[14]~FF  (.D(n950), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[14]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[14]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key1_counter[15]~FF  (.D(n955), .CE(n271), .CLK(\mipi_pclk~O ), 
           .SR(n874), .Q(\key1_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key1_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \key1_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \key1_counter[15]~FF .SR_POLARITY = 1'b1;
    defparam \key1_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \key1_counter[15]~FF .SR_SYNC = 1'b1;
    defparam \key1_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \key1_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[1]~FF  (.D(n379), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[1]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[1]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[1]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[1]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[1]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[1]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[2]~FF  (.D(n378), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[2]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[2]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[2]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[2]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[2]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[2]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[3]~FF  (.D(n377), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[3]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[3]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[3]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[3]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[3]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[3]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[4]~FF  (.D(n376), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[4]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[4]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[4]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[4]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[4]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[4]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[5]~FF  (.D(n375), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[5]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[5]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[5]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[5]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[5]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[5]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[6]~FF  (.D(n374), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[6]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[6]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[6]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[6]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[6]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[6]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[7]~FF  (.D(n373), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[7]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[7]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[7]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[7]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[7]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[7]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[8]~FF  (.D(n372), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[8]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[8]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[8]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[8]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[8]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[8]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[9]~FF  (.D(n371), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[9]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[9]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[9]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[9]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[9]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[9]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[10]~FF  (.D(n370), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[10]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[10]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[10]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[10]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[10]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[10]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[11]~FF  (.D(n369), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[11]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[11]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[11]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[11]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[11]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[11]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[12]~FF  (.D(n368), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[12]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[12]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[12]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[12]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[12]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[12]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[13]~FF  (.D(n367), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[13]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[13]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[13]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[13]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[13]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[13]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[14]~FF  (.D(n366), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[14]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[14]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[14]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[14]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[14]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[14]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \key2_counter[15]~FF  (.D(n365), .CE(ceg_net83), .CLK(\mipi_pclk~O ), 
           .SR(rx_status2), .Q(\key2_counter[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \key2_counter[15]~FF .CLK_POLARITY = 1'b1;
    defparam \key2_counter[15]~FF .CE_POLARITY = 1'b1;
    defparam \key2_counter[15]~FF .SR_POLARITY = 1'b0;
    defparam \key2_counter[15]~FF .D_POLARITY = 1'b1;
    defparam \key2_counter[15]~FF .SR_SYNC = 1'b1;
    defparam \key2_counter[15]~FF .SR_VALUE = 1'b0;
    defparam \key2_counter[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \red_gain[1]~FF  (.D(n390), .CE(\equal_59/n31 ), .CLK(\mipi_pclk~O ), 
           .SR(n875), .Q(\red_gain[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \red_gain[1]~FF .CLK_POLARITY = 1'b1;
    defparam \red_gain[1]~FF .CE_POLARITY = 1'b0;
    defparam \red_gain[1]~FF .SR_POLARITY = 1'b1;
    defparam \red_gain[1]~FF .D_POLARITY = 1'b1;
    defparam \red_gain[1]~FF .SR_SYNC = 1'b1;
    defparam \red_gain[1]~FF .SR_VALUE = 1'b0;
    defparam \red_gain[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \red_gain[2]~FF  (.D(n389), .CE(\equal_59/n31 ), .CLK(\mipi_pclk~O ), 
           .SR(n875), .Q(\red_gain[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b1, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \red_gain[2]~FF .CLK_POLARITY = 1'b1;
    defparam \red_gain[2]~FF .CE_POLARITY = 1'b0;
    defparam \red_gain[2]~FF .SR_POLARITY = 1'b1;
    defparam \red_gain[2]~FF .D_POLARITY = 1'b1;
    defparam \red_gain[2]~FF .SR_SYNC = 1'b1;
    defparam \red_gain[2]~FF .SR_VALUE = 1'b1;
    defparam \red_gain[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \green_gain[2]~FF  (.D(1'b1), .CE(n875), .CLK(\mipi_pclk~O ), 
           .SR(1'b0), .Q(\green_gain[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(199)
    defparam \green_gain[2]~FF .CLK_POLARITY = 1'b1;
    defparam \green_gain[2]~FF .CE_POLARITY = 1'b1;
    defparam \green_gain[2]~FF .SR_POLARITY = 1'b1;
    defparam \green_gain[2]~FF .D_POLARITY = 1'b1;
    defparam \green_gain[2]~FF .SR_SYNC = 1'b1;
    defparam \green_gain[2]~FF .SR_VALUE = 1'b0;
    defparam \green_gain[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[1]~FF  (.D(n141), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[1]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[1]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[2]~FF  (.D(n1062), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[2]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[2]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[3]~FF  (.D(n1060_2), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[3]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[3]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[4]~FF  (.D(n1058), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[4]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[4]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[5]~FF  (.D(n1056), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[5]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[6]~FF  (.D(n1028), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[6]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[7]~FF  (.D(n1026), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[7]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[8]~FF  (.D(n1000), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[8]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[8]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[9]~FF  (.D(n998), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[9]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[9]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[10]~FF  (.D(n995), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[10]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[10]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[10]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[10]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[10]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[10]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[11]~FF  (.D(n979), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[11]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[11]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[11]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[11]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[11]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[11]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_waddr_1P[12]~FF  (.D(n978), .CE(1'b1), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_waddr_1P[12]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_waddr_1P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \r_waddr_1P[12]~FF .CE_POLARITY = 1'b1;
    defparam \r_waddr_1P[12]~FF .SR_POLARITY = 1'b0;
    defparam \r_waddr_1P[12]~FF .D_POLARITY = 1'b1;
    defparam \r_waddr_1P[12]~FF .SR_SYNC = 1'b0;
    defparam \r_waddr_1P[12]~FF .SR_VALUE = 1'b0;
    defparam \r_waddr_1P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[0]~FF  (.D(\inst_line_buf/even_line_pix_0[0] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[0]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_valid_1P~FF  (.D(r_mipi_rx_valid_1P_2), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_valid_1P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_valid_1P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_valid_1P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_valid_1P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_valid_1P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_valid_1P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_valid_1P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_valid_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[0]~FF  (.D(\inst_line_buf/n1296 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[0]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[0]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[0]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[0]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[0]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_hsync_2P~FF  (.D(\inst_line_buf/r_mipi_rx_hsync_1P ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_hsync_2P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_hsync_2P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_hsync_2P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_hsync_2P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_hsync_2P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_hsync_2P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_hsync_2P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_hsync_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[0]~FF  (.D(\inst_line_buf/n1381 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[0]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[0]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[0]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_full_1P_2~FF  (.D(\inst_line_buf/r_mipi_rx_full_1P_2 ), 
           .CE(ceg_net101), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_full_1P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_full_1P_2~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_full_1P_2~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_full_1P_2~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_full_1P_2~FF .D_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_full_1P_2~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_full_1P_2~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_full_1P_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_en_1P~FF  (.D(\inst_line_buf/n2531 ), 
           .CE(ceg_net104), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_en_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_en_1P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_en_1P~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_en_1P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_en_1P~FF .D_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_en_1P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_en_1P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_en_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_inc_1P~FF  (.D(1'b1), .CE(\inst_line_buf/r_mipi_rx_full_1P_2 ), 
           .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_inc_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_inc_1P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_inc_1P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_inc_1P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_inc_1P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_inc_1P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_inc_1P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_inc_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_b_1P[0]~FF  (.D(\inst_line_buf/n1385 ), 
           .CE(ceg_net140), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_b_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_b_1P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_b_1P[0]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[0]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[0]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_b_1P[0]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[0]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[0]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[40] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[0]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[0]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[0]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[0]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[0]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[0]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_hsync_1P~FF  (.D(ceg_net140), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_hsync_1P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_hsync_1P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_1P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_1P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_1P~FF .D_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_1P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_1P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_valid_1P~FF  (.D(\inst_line_buf/n1387 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_valid_1P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_valid_1P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_1P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_1P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_1P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_1P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_1P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_hsync_2P~FF  (.D(\inst_line_buf/r_mipi_tx_hsync_1P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_hsync_2P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_hsync_2P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_2P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_2P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_2P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_2P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_2P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_valid_2P~FF  (.D(\inst_line_buf/r_mipi_tx_valid_1P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_valid_2P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_valid_2P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_2P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_2P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_2P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_2P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_2P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_2P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_hsync_3P~FF  (.D(\inst_line_buf/r_mipi_tx_hsync_2P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_hsync_3P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_hsync_3P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_3P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_3P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_3P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_3P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_3P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_3P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_valid_3P~FF  (.D(\inst_line_buf/r_mipi_tx_valid_2P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_valid_3P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_valid_3P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_3P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_3P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_3P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_3P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_3P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_3P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[0]~FF  (.D(\inst_line_buf/n1510 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[0])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[0]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[0]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[0]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[0]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[0]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[0]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[0]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_hsync_4P~FF  (.D(\inst_line_buf/r_mipi_tx_hsync_3P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_hsync_4P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_hsync_4P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_4P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_4P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_4P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_4P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_4P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_4P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_valid_4P~FF  (.D(\inst_line_buf/r_mipi_tx_valid_3P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_valid_4P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_valid_4P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_4P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_4P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_4P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_4P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_4P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_4P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_hsync_5P~FF  (.D(\inst_line_buf/r_mipi_tx_hsync_4P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_hsync_5P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_hsync_5P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_5P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_5P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_5P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_hsync_5P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_5P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_hsync_5P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_valid_5P~FF  (.D(\inst_line_buf/r_mipi_tx_valid_4P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_valid_5P_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_valid_5P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_5P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_5P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_5P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_valid_5P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_5P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_valid_5P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_hsync~FF  (.D(\inst_line_buf/r_mipi_tx_hsync_5P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(rx_status3)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_hsync~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_hsync~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_hsync~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_hsync~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_hsync~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_hsync~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_hsync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_valid~FF  (.D(\inst_line_buf/r_mipi_tx_valid_5P_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_VALID)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_valid~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_valid~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_valid~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_valid~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_valid~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_valid~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_valid~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_hsync_1P~FF  (.D(\r_mipi_rx_hsync_1P[0]_2 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_hsync_1P )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_hsync_1P~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_hsync_1P~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_hsync_1P~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_hsync_1P~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_hsync_1P~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_hsync_1P~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_hsync_1P~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[1]~FF  (.D(\inst_line_buf/odd_line_pix_0[1] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[1]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[1]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[2]~FF  (.D(\inst_line_buf/odd_line_pix_0[2] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[2]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[2]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[3]~FF  (.D(\inst_line_buf/odd_line_pix_0[3] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[3]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[3]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[4]~FF  (.D(\inst_line_buf/odd_line_pix_0[4] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[4]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[4]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[5]~FF  (.D(\inst_line_buf/odd_line_pix_0[5] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[5]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[5]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[6]~FF  (.D(\inst_line_buf/odd_line_pix_0[6] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[6]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[6]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[7]~FF  (.D(\inst_line_buf/odd_line_pix_0[7] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[7]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[7]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[8]~FF  (.D(\inst_line_buf/odd_line_pix_0[8] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[8]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[8]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[8]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[9]~FF  (.D(\inst_line_buf/odd_line_pix_0[9] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[9]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[9]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[9]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[10]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[10] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[10]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[10]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[10]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[10]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[10]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[10]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[11]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[11] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[11]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[11]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[11]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[11]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[11]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[11]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[12]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[12] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[12]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[12]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[12]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[12]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[12]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[12]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[13]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[13] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[13]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[13]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[13]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[13]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[13]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[13]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[13]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[14]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[14] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[14]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[14]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[14]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[14]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[14]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[14]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[14]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[15]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[15] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[15]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[15]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[15]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[15]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[15]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[15]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[15]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[16]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[16] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[16]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[16]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[16]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[16]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[16]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[16]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[16]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[17]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[17] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[17]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[17]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[17]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[17]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[17]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[17]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[17]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[18]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[18] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[18]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[18]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[18]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[18]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[18]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[18]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[18]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[19]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[19] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[19]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[19]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[19]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[19]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[19]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[19]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[19]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[20]~FF  (.D(\inst_line_buf/even_line_pix_2[0] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[20]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[20]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[20]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[20]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[20]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[20]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[20]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[21]~FF  (.D(\inst_line_buf/odd_line_pix_2[1] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[21]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[21]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[21]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[21]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[21]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[21]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[21]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[22]~FF  (.D(\inst_line_buf/odd_line_pix_2[2] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[22]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[22]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[22]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[22]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[22]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[22]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[22]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[23]~FF  (.D(\inst_line_buf/odd_line_pix_2[3] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[23]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[23]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[23]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[23]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[23]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[23]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[23]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[24]~FF  (.D(\inst_line_buf/odd_line_pix_2[4] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[24]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[24]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[24]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[24]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[24]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[24]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[24]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[25]~FF  (.D(\inst_line_buf/odd_line_pix_2[5] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[25]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[25]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[25]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[25]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[25]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[25]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[25]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[26]~FF  (.D(\inst_line_buf/odd_line_pix_2[6] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[26]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[26]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[26]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[26]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[26]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[26]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[26]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[27]~FF  (.D(\inst_line_buf/odd_line_pix_2[7] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[27]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[27]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[27]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[27]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[27]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[27]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[27]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[28]~FF  (.D(\inst_line_buf/odd_line_pix_2[8] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[28]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[28]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[28]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[28]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[28]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[28]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[28]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[29]~FF  (.D(\inst_line_buf/odd_line_pix_2[9] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[29]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[29]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[29]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[29]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[29]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[29]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[29]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[30]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[30] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[30]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[30]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[30]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[30]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[30]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[30]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[30]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[31]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[31] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[31]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[31]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[31]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[31]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[31]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[31]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[31]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[32]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[32] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[32]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[32]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[32]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[32]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[32]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[32]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[32]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[33]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[33] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[33]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[33]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[33]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[33]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[33]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[33]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[33]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[34]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[34] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[34]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[34]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[34]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[34]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[34]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[34]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[34]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[35]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[35] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[35]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[35]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[35]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[35]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[35]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[35]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[35]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[36]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[36] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[36]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[36]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[36]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[36]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[36]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[36]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[36]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[37]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[37] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[37]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[37]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[37]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[37]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[37]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[37]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[37]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[38]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[38] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[38]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[38]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[38]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[38]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[38]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[38]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[38]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_data_1P[39]~FF  (.D(\inst_line_buf/mipi_inst1_DATA_filtered[39] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_data_1P[39]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_data_1P[39]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[39]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[39]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[39]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_data_1P[39]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[39]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_data_1P[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[1]~FF  (.D(\inst_line_buf/n1295 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[1]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[1]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[1]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[1]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[1]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[1]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[2]~FF  (.D(\inst_line_buf/n1294 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[2]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[2]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[2]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[2]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[2]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[2]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[3]~FF  (.D(\inst_line_buf/n1293 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[3]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[3]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[3]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[3]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[3]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[3]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[4]~FF  (.D(\inst_line_buf/n1292 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[4]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[4]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[4]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[4]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[4]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[4]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[5]~FF  (.D(\inst_line_buf/n1291 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[5]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[5]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[5]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[5]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[5]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[5]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[6]~FF  (.D(\inst_line_buf/n1290 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[6]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[6]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[6]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[6]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[6]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[6]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[7]~FF  (.D(\inst_line_buf/n1289 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[7]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[7]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[7]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[7]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[7]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[7]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[8]~FF  (.D(\inst_line_buf/n1288 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[8]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[8]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[8]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[8]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[8]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[8]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[9]~FF  (.D(\inst_line_buf/n1287 ), 
           .CE(ceg_net98), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_rx_x_2P[9]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[9]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[9]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[9]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[9]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[9]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF  (.D(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
           .CE(\inst_line_buf/n1283 ), .CLK(\mipi_pclk~O ), .SR(rx_status2), 
           .Q(\inst_line_buf/r_mipi_rx_x_2P[10]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF .D_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_rx_x_2P[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[1]~FF  (.D(\inst_line_buf/n1380 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[1]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[1]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[2]~FF  (.D(\inst_line_buf/n1379 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[2]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[2]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[3]~FF  (.D(\inst_line_buf/n1378 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[3]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[3]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[4]~FF  (.D(\inst_line_buf/n1377 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[4]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[4]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[5]~FF  (.D(\inst_line_buf/n1376 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[5]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[5]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[6]~FF  (.D(\inst_line_buf/n1375 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[6]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[6]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[7]~FF  (.D(\inst_line_buf/n1374 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[7]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[7]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[8]~FF  (.D(\inst_line_buf/n1373 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[8]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[8]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[8]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[9]~FF  (.D(\inst_line_buf/n1372 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_x_1P[9]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[9]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[9]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF  (.D(\inst_line_buf/r_mipi_tx_x_1P[10]_2 ), 
           .CE(\inst_line_buf/n2531 ), .CLK(\mipi_pclk~O ), .SR(rx_status2), 
           .Q(\inst_line_buf/r_mipi_tx_x_1P[10]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b0, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF .D_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_x_1P[10]_2~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_b_1P[1]~FF  (.D(\inst_line_buf/n1384 ), 
           .CE(ceg_net140), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_b_1P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_b_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_b_1P[1]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[1]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_b_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_b_1P[2]~FF  (.D(\inst_line_buf/n1383 ), 
           .CE(ceg_net140), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_b_1P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b0, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_b_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_b_1P[2]~FF .CE_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[2]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_b_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_b_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[1]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[41] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[1]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[1]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[1]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[1]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[1]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[2]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[42] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[2]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[2]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[2]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[2]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[2]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[3]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[43] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[3]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[3]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[3]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[3]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[3]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[4]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[44] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[4]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[4]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[4]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[4]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[4]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[5]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[45] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[5]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[5]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[5]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[5]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[5]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[6]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[46] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[6]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[6]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[6]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[6]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[6]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[7]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[47] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[7]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[7]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[7]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[7]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[7]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[8]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[48] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[8]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[8]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[8]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[8]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[8]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[9]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[49] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[9]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[9]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[9]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[9]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[9]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[10]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[50] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[10]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[10]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[10]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[10]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[10]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[11]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[51] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[11]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[11]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[11]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[11]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[11]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[12]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[52] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[12]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[12]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[12]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[12]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[12]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[13]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[53] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[13]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[13]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[13]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[13]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[13]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[13]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[14]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[54] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[14]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[14]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[14]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[14]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[14]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[14]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[15]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[55] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[15]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[15]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[15]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[15]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[15]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[15]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[16]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[56] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[16]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[16]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[16]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[16]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[16]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[16]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[17]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[57] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[17]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[17]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[17]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[17]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[17]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[17]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[18]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[58] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[18]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[18]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[18]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[18]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[18]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[18]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[19]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[59] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[19]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[19]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[19]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[19]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[19]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[19]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[20]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[60] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[20] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[20]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[20]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[20]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[20]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[20]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[20]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[21]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[61] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[21] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[21]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[21]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[21]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[21]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[21]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[21]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[22]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[62] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[22] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[22]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[22]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[22]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[22]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[22]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[22]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[23]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[63] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[23] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[23]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[23]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[23]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[23]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[23]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[23]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[24]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[64] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[24] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[24]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[24]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[24]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[24]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[24]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[24]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[25]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[65] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[25] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[25]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[25]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[25]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[25]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[25]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[25]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[26]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[66] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[26] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[26]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[26]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[26]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[26]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[26]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[26]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[27]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[67] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[27] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[27]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[27]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[27]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[27]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[27]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[27]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[28]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[68] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[28] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[28]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[28]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[28]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[28]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[28]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[28]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[29]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[69] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[29] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[29]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[29]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[29]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[29]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[29]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[29]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[30]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[70] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[30]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[30]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[30]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[30]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[30]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[30]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[31]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[71] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[31]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[31]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[31]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[31]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[31]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[31]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[32]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[72] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[32]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[32]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[32]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[32]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[32]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[32]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[33]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[73] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[33]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[33]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[33]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[33]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[33]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[33]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[34]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[74] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[34]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[34]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[34]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[34]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[34]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[34]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[35]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[75] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[35]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[35]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[35]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[35]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[35]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[35]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[36]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[76] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[36]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[36]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[36]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[36]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[36]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[36]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[37]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[77] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[37]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[37]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[37]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[37]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[37]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[37]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[38]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[78] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[38]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[38]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[38]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[38]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[38]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[38]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[39]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[79] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[39]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[39]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[39]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[39]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[39]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[39]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[40]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[80] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[40] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[40]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[40]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[40]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[40]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[40]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[40]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[41]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[81] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[41] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[41]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[41]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[41]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[41]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[41]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[41]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[42]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[82] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[42] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[42]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[42]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[42]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[42]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[42]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[42]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[43]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[83] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[43] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[43]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[43]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[43]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[43]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[43]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[43]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[44]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[84] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[44] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[44]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[44]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[44]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[44]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[44]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[44]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[45]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[85] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[45] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[45]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[45]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[45]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[45]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[45]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[45]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[46]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[86] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[46] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[46]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[46]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[46]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[46]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[46]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[46]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[47]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[87] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[47] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[47]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[47]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[47]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[47]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[47]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[47]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[48]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[88] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[48] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[48]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[48]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[48]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[48]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[48]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[48]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[49]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[89] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[49] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[49]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[49]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[49]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[49]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[49]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[49]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[50]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[90] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[50] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[50]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[50]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[50]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[50]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[50]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[50]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[51]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[91] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[51] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[51]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[51]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[51]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[51]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[51]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[51]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[52]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[92] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[52] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[52]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[52]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[52]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[52]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[52]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[52]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[53]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[93] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[53] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[53]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[53]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[53]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[53]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[53]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[53]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[54]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[94] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[54] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[54]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[54]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[54]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[54]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[54]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[54]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[55]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[95] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[55] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[55]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[55]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[55]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[55]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[55]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[55]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[56]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[96] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[56] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[56]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[56]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[56]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[56]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[56]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[56]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[57]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[97] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[57] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[57]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[57]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[57]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[57]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[57]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[57]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[58]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[98] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[58] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[58]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[58]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[58]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[58]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[58]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[58]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[59]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[99] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[59] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[59]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[59]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[59]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[59]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[59]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[59]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[60]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[100] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[60]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[60]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[60]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[60]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[60]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[60]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[61]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[101] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[61]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[61]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[61]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[61]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[61]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[61]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[62]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[102] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[62]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[62]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[62]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[62]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[62]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[62]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[63]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[103] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[63]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[63]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[63]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[63]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[63]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[63]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[64]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[104] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[64]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[64]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[64]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[64]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[64]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[64]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[65]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[105] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[65]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[65]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[65]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[65]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[65]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[65]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[66]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[106] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[66]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[66]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[66]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[66]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[66]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[66]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[67]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[107] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[67]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[67]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[67]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[67]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[67]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[67]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[68]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[108] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[68]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[68]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[68]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[68]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[68]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[68]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[69]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[109] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[69]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[69]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[69]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[69]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[69]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[69]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[70]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[110] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[70]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[70]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[70]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[70]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[70]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[70]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[71]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[111] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[71]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[71]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[71]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[71]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[71]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[71]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[72]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[112] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[72]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[72]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[72]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[72]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[72]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[72]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[73]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[113] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[73]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[73]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[73]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[73]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[73]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[73]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[74]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[114] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[74]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[74]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[74]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[74]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[74]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[74]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[75]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[115] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[75]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[75]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[75]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[75]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[75]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[75]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[76]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[116] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[76]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[76]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[76]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[76]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[76]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[76]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[77]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[117] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[77]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[77]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[77]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[77]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[77]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[77]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[78]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[118] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[78]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[78]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[78]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[78]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[78]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[78]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[79]~FF  (.D(\inst_line_buf/r_mipi_tx_data_4P[119] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[79]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[79]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[79]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[79]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[79]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[79]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[80]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[0] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[80]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[80]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[80]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[80]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[80]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[80]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[81]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[1] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[81]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[81]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[81]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[81]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[81]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[81]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[82]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[2] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[82]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[82]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[82]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[82]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[82]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[82]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[83]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[3] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[83]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[83]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[83]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[83]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[83]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[83]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[84]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[4] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[84]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[84]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[84]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[84]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[84]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[84]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[85]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[5] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[85]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[85]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[85]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[85]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[85]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[85]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[86]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[6] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[86]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[86]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[86]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[86]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[86]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[86]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[87]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[7] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[87]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[87]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[87]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[87]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[87]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[87]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[88]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[8] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[88]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[88]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[88]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[88]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[88]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[88]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[89]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[9] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[89]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[89]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[89]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[89]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[89]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[89]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[90]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[10] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[90]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[90]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[90]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[90]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[90]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[90]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[91]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[11] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[91]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[91]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[91]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[91]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[91]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[91]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[92]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[12] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[92]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[92]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[92]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[92]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[92]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[92]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[93]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[13] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[93]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[93]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[93]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[93]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[93]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[93]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[94]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[14] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[94]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[94]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[94]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[94]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[94]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[94]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[95]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[15] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[95]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[95]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[95]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[95]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[95]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[95]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[96]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[16] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[96]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[96]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[96]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[96]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[96]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[96]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[97]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[17] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[97]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[97]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[97]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[97]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[97]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[97]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[98]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[18] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[98]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[98]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[98]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[98]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[98]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[98]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[99]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[19] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[99]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[99]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[99]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[99]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[99]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[99]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[100]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[20] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[100]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[100]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[100]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[100]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[100]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[100]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[101]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[21] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[101]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[101]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[101]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[101]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[101]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[101]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[102]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[22] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[102]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[102]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[102]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[102]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[102]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[102]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[103]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[23] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[103]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[103]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[103]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[103]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[103]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[103]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[104]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[24] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[104]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[104]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[104]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[104]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[104]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[104]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[105]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[25] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[105]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[105]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[105]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[105]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[105]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[105]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[106]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[26] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[106]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[106]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[106]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[106]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[106]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[106]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[107]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[27] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[107]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[107]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[107]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[107]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[107]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[107]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[108]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[28] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[108]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[108]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[108]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[108]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[108]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[108]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[109]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[29] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[109]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[109]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[109]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[109]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[109]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[109]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[110]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[30] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[110]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[110]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[110]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[110]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[110]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[110]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[111]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[31] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[111]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[111]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[111]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[111]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[111]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[111]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[112]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[32] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[112]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[112]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[112]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[112]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[112]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[112]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[113]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[33] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[113]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[113]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[113]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[113]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[113]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[113]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[114]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[34] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[114]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[114]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[114]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[114]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[114]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[114]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[115]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[35] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[115]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[115]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[115]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[115]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[115]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[115]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[116]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[36] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[116]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[116]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[116]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[116]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[116]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[116]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[117]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[37] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[117]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[117]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[117]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[117]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[117]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[117]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[118]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[38] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[118]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[118]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[118]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[118]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[118]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[118]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_4P[119]~FF  (.D(\inst_line_buf/w_mipi_tx_data_3P[39] ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_4P[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_4P[119]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[119]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[119]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[119]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_4P[119]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[119]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_4P[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[1]~FF  (.D(\inst_line_buf/n1509 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[1])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[1]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[1]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[1]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[1]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[1]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[1]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[2]~FF  (.D(\inst_line_buf/n1508 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[2])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[2]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[2]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[2]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[2]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[2]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[2]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[3]~FF  (.D(\inst_line_buf/n1507 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[3])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[3]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[3]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[3]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[3]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[3]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[3]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[4]~FF  (.D(\inst_line_buf/n1506 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[4])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[4]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[4]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[4]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[4]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[4]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[4]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[5]~FF  (.D(\inst_line_buf/n1505 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[5])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[5]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[5]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[5]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[5]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[5]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[5]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[6]~FF  (.D(\inst_line_buf/n1504 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[6])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[6]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[6]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[6]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[6]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[6]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[6]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[7]~FF  (.D(\inst_line_buf/n1503 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[7])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[7]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[7]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[7]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[7]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[7]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[7]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[8]~FF  (.D(\inst_line_buf/n1502 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[8])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[8]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[8]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[8]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[8]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[8]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[8]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[9]~FF  (.D(\inst_line_buf/n1501 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[9])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[9]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[9]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[9]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[9]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[9]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[9]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[10]~FF  (.D(\inst_line_buf/n1500 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[10])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[10]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[10]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[10]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[10]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[10]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[10]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[11]~FF  (.D(\inst_line_buf/n1499 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[11])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[11]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[11]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[11]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[11]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[11]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[11]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[12]~FF  (.D(\inst_line_buf/n1498 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[12])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[12]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[12]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[12]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[12]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[12]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[12]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[13]~FF  (.D(\inst_line_buf/n1497 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[13])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[13]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[13]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[13]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[13]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[13]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[13]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[13]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[14]~FF  (.D(\inst_line_buf/n1496 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[14])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[14]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[14]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[14]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[14]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[14]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[14]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[14]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[15]~FF  (.D(\inst_line_buf/n1495 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[15])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[15]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[15]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[15]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[15]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[15]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[15]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[15]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[16]~FF  (.D(\inst_line_buf/n1494 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[16])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[16]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[16]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[16]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[16]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[16]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[16]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[16]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[17]~FF  (.D(\inst_line_buf/n1493 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[17])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[17]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[17]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[17]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[17]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[17]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[17]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[17]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[18]~FF  (.D(\inst_line_buf/n1492 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[18])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[18]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[18]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[18]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[18]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[18]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[18]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[18]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[19]~FF  (.D(\inst_line_buf/n1491 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[19])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[19]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[19]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[19]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[19]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[19]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[19]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[19]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[20]~FF  (.D(\inst_line_buf/n1490 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[20])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[20]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[20]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[20]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[20]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[20]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[20]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[20]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[21]~FF  (.D(\inst_line_buf/n1489 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[21])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[21]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[21]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[21]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[21]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[21]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[21]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[21]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[22]~FF  (.D(\inst_line_buf/n1488 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[22])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[22]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[22]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[22]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[22]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[22]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[22]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[22]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[23]~FF  (.D(\inst_line_buf/n1487 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[23])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[23]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[23]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[23]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[23]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[23]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[23]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[23]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[24]~FF  (.D(\inst_line_buf/n1486 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[24])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[24]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[24]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[24]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[24]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[24]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[24]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[24]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[25]~FF  (.D(\inst_line_buf/n1485 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[25])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[25]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[25]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[25]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[25]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[25]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[25]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[25]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[26]~FF  (.D(\inst_line_buf/n1484 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[26])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[26]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[26]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[26]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[26]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[26]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[26]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[26]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[27]~FF  (.D(\inst_line_buf/n1483 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[27])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[27]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[27]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[27]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[27]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[27]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[27]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[27]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[28]~FF  (.D(\inst_line_buf/n1482 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[28])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[28]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[28]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[28]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[28]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[28]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[28]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[28]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[29]~FF  (.D(\inst_line_buf/n1481 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[29])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[29]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[29]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[29]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[29]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[29]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[29]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[29]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[30]~FF  (.D(\inst_line_buf/n1480 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[30])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[30]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[30]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[30]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[30]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[30]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[30]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[30]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[31]~FF  (.D(\inst_line_buf/n1479 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[31])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[31]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[31]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[31]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[31]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[31]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[31]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[31]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[32]~FF  (.D(\inst_line_buf/n1478 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[32])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[32]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[32]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[32]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[32]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[32]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[32]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[32]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[33]~FF  (.D(\inst_line_buf/n1477 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[33])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[33]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[33]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[33]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[33]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[33]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[33]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[33]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[34]~FF  (.D(\inst_line_buf/n1476 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[34])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[34]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[34]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[34]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[34]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[34]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[34]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[34]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[35]~FF  (.D(\inst_line_buf/n1475 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[35])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[35]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[35]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[35]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[35]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[35]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[35]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[35]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[36]~FF  (.D(\inst_line_buf/n1474 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[36])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[36]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[36]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[36]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[36]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[36]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[36]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[36]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[37]~FF  (.D(\inst_line_buf/n1473 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[37])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[37]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[37]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[37]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[37]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[37]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[37]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[37]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[38]~FF  (.D(\inst_line_buf/n1472 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[38])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[38]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[38]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[38]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[38]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[38]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[38]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[38]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[39]~FF  (.D(\inst_line_buf/n1471 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[39])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[39]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[39]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[39]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[39]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[39]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[39]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[39]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[40]~FF  (.D(\inst_line_buf/n1470 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[40])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[40]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[40]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[40]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[40]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[40]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[40]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[40]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[41]~FF  (.D(\inst_line_buf/n1469 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[41])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[41]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[41]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[41]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[41]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[41]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[41]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[41]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[42]~FF  (.D(\inst_line_buf/n1468 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[42])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[42]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[42]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[42]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[42]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[42]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[42]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[42]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[43]~FF  (.D(\inst_line_buf/n1467 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[43])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[43]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[43]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[43]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[43]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[43]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[43]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[43]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[44]~FF  (.D(\inst_line_buf/n1466 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[44])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[44]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[44]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[44]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[44]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[44]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[44]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[44]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[45]~FF  (.D(\inst_line_buf/n1465 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[45])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[45]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[45]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[45]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[45]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[45]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[45]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[45]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[46]~FF  (.D(\inst_line_buf/n1464 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[46])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[46]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[46]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[46]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[46]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[46]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[46]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[46]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[47]~FF  (.D(\inst_line_buf/n1463 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[47])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[47]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[47]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[47]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[47]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[47]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[47]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[47]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[48]~FF  (.D(\inst_line_buf/n1462 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[48])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[48]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[48]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[48]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[48]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[48]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[48]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[48]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[49]~FF  (.D(\inst_line_buf/n1461 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[49])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[49]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[49]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[49]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[49]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[49]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[49]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[49]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[50]~FF  (.D(\inst_line_buf/n1460 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[50])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[50]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[50]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[50]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[50]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[50]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[50]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[50]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[51]~FF  (.D(\inst_line_buf/n1459 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[51])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[51]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[51]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[51]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[51]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[51]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[51]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[51]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[52]~FF  (.D(\inst_line_buf/n1458 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[52])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[52]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[52]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[52]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[52]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[52]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[52]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[52]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[53]~FF  (.D(\inst_line_buf/n1457 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[53])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[53]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[53]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[53]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[53]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[53]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[53]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[53]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[54]~FF  (.D(\inst_line_buf/n1456 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[54])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[54]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[54]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[54]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[54]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[54]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[54]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[54]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[55]~FF  (.D(\inst_line_buf/n1455 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[55])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[55]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[55]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[55]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[55]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[55]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[55]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[55]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[56]~FF  (.D(\inst_line_buf/n1454 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[56])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[56]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[56]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[56]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[56]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[56]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[56]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[56]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[57]~FF  (.D(\inst_line_buf/n1453 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[57])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[57]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[57]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[57]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[57]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[57]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[57]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[57]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[58]~FF  (.D(\inst_line_buf/n1452 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[58])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[58]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[58]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[58]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[58]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[58]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[58]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[58]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/w_mipi_tx_data[59]~FF  (.D(\inst_line_buf/n1451 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(mipi_inst2_DATA[59])) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/w_mipi_tx_data[59]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[59]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[59]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[59]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/w_mipi_tx_data[59]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[59]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/w_mipi_tx_data[59]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[60]~FF  (.D(\inst_line_buf/n1450 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[60] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[60]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[60]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[60]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[60]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[60]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[60]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[60]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[61]~FF  (.D(\inst_line_buf/n1449 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[61] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[61]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[61]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[61]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[61]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[61]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[61]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[61]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[62]~FF  (.D(\inst_line_buf/n1448 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[62] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[62]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[62]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[62]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[62]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[62]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[62]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[62]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[63]~FF  (.D(\inst_line_buf/n1447 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[63] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[63]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[63]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[63]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[63]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[63]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[63]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[63]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[64]~FF  (.D(\inst_line_buf/n1446 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[64] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[64]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[64]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[64]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[64]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[64]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[64]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[64]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[65]~FF  (.D(\inst_line_buf/n1445 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[65] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[65]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[65]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[65]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[65]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[65]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[65]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[65]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[66]~FF  (.D(\inst_line_buf/n1444 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[66] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[66]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[66]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[66]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[66]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[66]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[66]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[66]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[67]~FF  (.D(\inst_line_buf/n1443 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[67] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[67]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[67]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[67]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[67]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[67]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[67]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[67]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[68]~FF  (.D(\inst_line_buf/n1442 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[68] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[68]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[68]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[68]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[68]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[68]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[68]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[68]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[69]~FF  (.D(\inst_line_buf/n1441 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[69] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[69]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[69]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[69]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[69]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[69]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[69]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[69]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[70]~FF  (.D(\inst_line_buf/n1440 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[70] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[70]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[70]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[70]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[70]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[70]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[70]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[70]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[71]~FF  (.D(\inst_line_buf/n1439 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[71] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[71]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[71]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[71]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[71]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[71]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[71]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[71]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[72]~FF  (.D(\inst_line_buf/n1438 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[72] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[72]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[72]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[72]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[72]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[72]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[72]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[72]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[73]~FF  (.D(\inst_line_buf/n1437 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[73] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[73]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[73]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[73]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[73]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[73]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[73]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[73]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[74]~FF  (.D(\inst_line_buf/n1436 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[74] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[74]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[74]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[74]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[74]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[74]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[74]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[74]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[75]~FF  (.D(\inst_line_buf/n1435 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[75] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[75]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[75]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[75]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[75]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[75]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[75]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[75]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[76]~FF  (.D(\inst_line_buf/n1434 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[76] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[76]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[76]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[76]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[76]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[76]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[76]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[76]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[77]~FF  (.D(\inst_line_buf/n1433 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[77] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[77]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[77]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[77]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[77]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[77]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[77]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[77]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[78]~FF  (.D(\inst_line_buf/n1432 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[78] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[78]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[78]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[78]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[78]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[78]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[78]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[78]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[79]~FF  (.D(\inst_line_buf/n1431 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[79] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[79]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[79]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[79]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[79]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[79]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[79]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[79]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[80]~FF  (.D(\inst_line_buf/n1430 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[80] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[80]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[80]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[80]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[80]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[80]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[80]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[80]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[81]~FF  (.D(\inst_line_buf/n1429 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[81] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[81]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[81]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[81]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[81]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[81]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[81]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[81]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[82]~FF  (.D(\inst_line_buf/n1428 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[82] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[82]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[82]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[82]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[82]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[82]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[82]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[82]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[83]~FF  (.D(\inst_line_buf/n1427 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[83] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[83]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[83]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[83]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[83]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[83]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[83]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[83]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[84]~FF  (.D(\inst_line_buf/n1426 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[84] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[84]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[84]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[84]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[84]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[84]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[84]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[84]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[85]~FF  (.D(\inst_line_buf/n1425 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[85] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[85]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[85]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[85]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[85]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[85]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[85]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[85]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[86]~FF  (.D(\inst_line_buf/n1424 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[86] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[86]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[86]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[86]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[86]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[86]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[86]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[86]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[87]~FF  (.D(\inst_line_buf/n1423 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[87] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[87]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[87]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[87]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[87]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[87]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[87]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[87]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[88]~FF  (.D(\inst_line_buf/n1422 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[88] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[88]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[88]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[88]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[88]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[88]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[88]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[88]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[89]~FF  (.D(\inst_line_buf/n1421 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[89] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[89]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[89]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[89]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[89]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[89]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[89]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[89]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[90]~FF  (.D(\inst_line_buf/n1420 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[90] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[90]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[90]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[90]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[90]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[90]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[90]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[90]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[91]~FF  (.D(\inst_line_buf/n1419 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[91] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[91]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[91]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[91]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[91]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[91]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[91]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[91]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[92]~FF  (.D(\inst_line_buf/n1418 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[92] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[92]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[92]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[92]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[92]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[92]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[92]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[92]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[93]~FF  (.D(\inst_line_buf/n1417 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[93] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[93]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[93]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[93]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[93]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[93]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[93]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[93]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[94]~FF  (.D(\inst_line_buf/n1416 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[94] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[94]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[94]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[94]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[94]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[94]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[94]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[94]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[95]~FF  (.D(\inst_line_buf/n1415 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[95] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[95]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[95]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[95]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[95]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[95]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[95]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[95]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[96]~FF  (.D(\inst_line_buf/n1414 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[96] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[96]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[96]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[96]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[96]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[96]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[96]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[96]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[97]~FF  (.D(\inst_line_buf/n1413 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[97] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[97]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[97]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[97]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[97]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[97]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[97]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[97]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[98]~FF  (.D(\inst_line_buf/n1412 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[98] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[98]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[98]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[98]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[98]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[98]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[98]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[98]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[99]~FF  (.D(\inst_line_buf/n1411 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[99] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[99]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[99]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[99]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[99]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[99]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[99]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[99]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[100]~FF  (.D(\inst_line_buf/n1410 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[100] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[100]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[100]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[100]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[100]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[100]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[100]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[100]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[101]~FF  (.D(\inst_line_buf/n1409 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[101] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[101]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[101]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[101]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[101]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[101]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[101]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[101]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[102]~FF  (.D(\inst_line_buf/n1408 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[102] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[102]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[102]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[102]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[102]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[102]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[102]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[102]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[103]~FF  (.D(\inst_line_buf/n1407 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[103] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[103]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[103]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[103]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[103]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[103]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[103]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[103]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[104]~FF  (.D(\inst_line_buf/n1406 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[104] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[104]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[104]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[104]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[104]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[104]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[104]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[104]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[105]~FF  (.D(\inst_line_buf/n1405 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[105] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[105]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[105]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[105]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[105]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[105]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[105]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[105]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[106]~FF  (.D(\inst_line_buf/n1404 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[106] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[106]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[106]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[106]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[106]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[106]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[106]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[106]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[107]~FF  (.D(\inst_line_buf/n1403 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[107] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[107]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[107]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[107]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[107]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[107]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[107]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[107]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[108]~FF  (.D(\inst_line_buf/n1402 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[108] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[108]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[108]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[108]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[108]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[108]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[108]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[108]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[109]~FF  (.D(\inst_line_buf/n1401 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[109] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[109]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[109]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[109]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[109]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[109]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[109]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[109]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[110]~FF  (.D(\inst_line_buf/n1400 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[110] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[110]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[110]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[110]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[110]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[110]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[110]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[110]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[111]~FF  (.D(\inst_line_buf/n1399 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[111] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[111]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[111]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[111]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[111]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[111]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[111]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[111]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[112]~FF  (.D(\inst_line_buf/n1398 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[112] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[112]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[112]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[112]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[112]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[112]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[112]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[112]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[113]~FF  (.D(\inst_line_buf/n1397 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[113] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[113]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[113]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[113]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[113]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[113]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[113]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[113]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[114]~FF  (.D(\inst_line_buf/n1396 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[114] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[114]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[114]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[114]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[114]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[114]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[114]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[114]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[115]~FF  (.D(\inst_line_buf/n1395 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[115] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[115]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[115]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[115]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[115]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[115]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[115]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[115]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[116]~FF  (.D(\inst_line_buf/n1394 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[116] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[116]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[116]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[116]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[116]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[116]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[116]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[116]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[117]~FF  (.D(\inst_line_buf/n1393 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[117] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[117]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[117]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[117]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[117]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[117]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[117]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[117]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[118]~FF  (.D(\inst_line_buf/n1392 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[118] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[118]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[118]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[118]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[118]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[118]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[118]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[118]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_line_buf/r_mipi_tx_data_5P[119]~FF  (.D(\inst_line_buf/n1391 ), 
           .CE(1'b1), .CLK(\mipi_pclk~O ), .SR(rx_status2), .Q(\inst_line_buf/r_mipi_tx_data_5P[119] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(296)
    defparam \inst_line_buf/r_mipi_tx_data_5P[119]~FF .CLK_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[119]~FF .CE_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[119]~FF .SR_POLARITY = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[119]~FF .D_POLARITY = 1'b1;
    defparam \inst_line_buf/r_mipi_tx_data_5P[119]~FF .SR_SYNC = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[119]~FF .SR_VALUE = 1'b0;
    defparam \inst_line_buf/r_mipi_tx_data_5P[119]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_GBUFCE CLKBUF__0 (.CE(1'b1), .I(mipi_pclk), .O(\mipi_pclk~O )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_GBUFCE, CE_POLARITY=1'b1 */ ;
    defparam CLKBUF__0.CE_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__inst_line_buf/add_64/i10  (.I0(1'b0), .I1(1'b0), 
            .CI(n2442), .O(n961)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \AUX_ADD_CO__inst_line_buf/add_64/i10 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__inst_line_buf/add_64/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CO__inst_line_buf/add_88/i10  (.I0(1'b0), .I1(1'b0), 
            .CI(n2441), .O(n903)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \AUX_ADD_CO__inst_line_buf/add_88/i10 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CO__inst_line_buf/add_88/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_97/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2440)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \AUX_ADD_CI__inst_line_buf/sub_97/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_97/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_94/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2439)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \AUX_ADD_CI__inst_line_buf/sub_94/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_94/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_82/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2438)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \AUX_ADD_CI__inst_line_buf/sub_82/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_82/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_73/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2437)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \AUX_ADD_CI__inst_line_buf/sub_73/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_73/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_70/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2436)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \AUX_ADD_CI__inst_line_buf/sub_70/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_70/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_61/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2435)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \AUX_ADD_CI__inst_line_buf/sub_61/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_61/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_58/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2434)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \AUX_ADD_CI__inst_line_buf/sub_58/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_58/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_55/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2433)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \AUX_ADD_CI__inst_line_buf/sub_55/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_55/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_49/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2432)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \AUX_ADD_CI__inst_line_buf/sub_49/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_49/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_46/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2431)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \AUX_ADD_CI__inst_line_buf/sub_46/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_46/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_43/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2430)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \AUX_ADD_CI__inst_line_buf/sub_43/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_43/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_37/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2429)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \AUX_ADD_CI__inst_line_buf/sub_37/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_37/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_31/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2428)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \AUX_ADD_CI__inst_line_buf/sub_31/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_31/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_22/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2427)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \AUX_ADD_CI__inst_line_buf/sub_22/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_22/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_25/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2426)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \AUX_ADD_CI__inst_line_buf/sub_25/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_25/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \AUX_ADD_CI__inst_line_buf/sub_19/add_2/i1  (.I0(1'b1), .I1(1'b1), 
            .CI(1'b0), .CO(n2425)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \AUX_ADD_CI__inst_line_buf/sub_19/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \AUX_ADD_CI__inst_line_buf/sub_19/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_FF \r_raddr_1P[1]~FF  (.D(n1060), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[1]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[1]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[1]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[1]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[1]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[1]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[1]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[1]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[2]~FF  (.D(n1065), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[2]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[2]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[2]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[2]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[2]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[2]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[2]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[2]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[3]~FF  (.D(n1070), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[3]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[3]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[3]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[3]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[3]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[3]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[3]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[3]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[4]~FF  (.D(n1075), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[4]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[4]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[4]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[4]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[4]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[4]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[4]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[4]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[5]~FF  (.D(n1080), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[5]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[5]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[5]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[5]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[5]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[5]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[5]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[5]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[6]~FF  (.D(n1085), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[6]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[6]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[6]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[6]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[6]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[6]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[6]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[6]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[7]~FF  (.D(n1090), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[7]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[7]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[7]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[7]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[7]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[7]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[7]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[7]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[8]~FF  (.D(n1095), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[8]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[8]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[8]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[8]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[8]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[8]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[8]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[8]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[9]~FF  (.D(n1100), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[9]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[9]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[9]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[9]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[9]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[9]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[9]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[9]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[10]~FF  (.D(n1105), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[10]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[10]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[10]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[10]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[10]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[10]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[10]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[10]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[11]~FF  (.D(n1110), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[11]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[11]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[11]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[11]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[11]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[11]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[11]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[11]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \r_raddr_1P[12]~FF  (.D(n1115), .CE(r_rden_1P_2), .CLK(\mipi_pclk~O ), 
           .SR(i_arstn), .Q(\r_raddr_1P[12]_2 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b0, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(249)
    defparam \r_raddr_1P[12]~FF .CLK_POLARITY = 1'b1;
    defparam \r_raddr_1P[12]~FF .CE_POLARITY = 1'b1;
    defparam \r_raddr_1P[12]~FF .SR_POLARITY = 1'b0;
    defparam \r_raddr_1P[12]~FF .D_POLARITY = 1'b1;
    defparam \r_raddr_1P[12]~FF .SR_SYNC = 1'b0;
    defparam \r_raddr_1P[12]~FF .SR_VALUE = 1'b0;
    defparam \r_raddr_1P[12]~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_dly/w_mipi_tx_vsync~FF  (.D(\inst_dly/r_rdata_1P[0] ), .CE(1'b1), 
           .CLK(\mipi_pclk~O ), .SR(1'b0), .Q(mipi_inst2_VSYNC)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(54)
    defparam \inst_dly/w_mipi_tx_vsync~FF .CLK_POLARITY = 1'b1;
    defparam \inst_dly/w_mipi_tx_vsync~FF .CE_POLARITY = 1'b1;
    defparam \inst_dly/w_mipi_tx_vsync~FF .SR_POLARITY = 1'b1;
    defparam \inst_dly/w_mipi_tx_vsync~FF .D_POLARITY = 1'b1;
    defparam \inst_dly/w_mipi_tx_vsync~FF .SR_SYNC = 1'b1;
    defparam \inst_dly/w_mipi_tx_vsync~FF .SR_VALUE = 1'b0;
    defparam \inst_dly/w_mipi_tx_vsync~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_FF \inst_dly/n24~FF  (.D(\r_raddr_1P[12]_2 ), .CE(r_rden_1P_2), 
           .CLK(\mipi_pclk~O ), .SR(1'b0), .Q(\inst_dly/n24 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_FF, CLK_POLARITY=1'b1, D_POLARITY=1'b1, CE_POLARITY=1'b1, SR_SYNC=1'b1, SR_SYNC_PRIORITY=1'b1, SR_VALUE=1'b0, SR_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(52)
    defparam \inst_dly/n24~FF .CLK_POLARITY = 1'b1;
    defparam \inst_dly/n24~FF .CE_POLARITY = 1'b1;
    defparam \inst_dly/n24~FF .SR_POLARITY = 1'b1;
    defparam \inst_dly/n24~FF .D_POLARITY = 1'b1;
    defparam \inst_dly/n24~FF .SR_SYNC = 1'b1;
    defparam \inst_dly/n24~FF .SR_VALUE = 1'b0;
    defparam \inst_dly/n24~FF .SR_SYNC_PRIORITY = 1'b1;
    EFX_ADD \add_81/i2  (.I0(\r_waddr_1P[1]_2 ), .I1(\r_waddr_1P[0]_2 ), 
            .CI(1'b0), .O(n141), .CO(n142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i2 .I0_POLARITY = 1'b1;
    defparam \add_81/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i4  (.I0(n200), .I1(n1247), .CI(n154), 
            .O(n150), .CO(n151)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i3  (.I0(n202), .I1(n1251), .CI(n156), 
            .O(n153), .CO(n154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i2  (.I0(n204), .I1(n1254), .CI(n418), 
            .O(n155), .CO(n156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i11  (.I0(n864), .I1(1'b1), .CI(n159_2), 
            .O(n157)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i10  (.I0(n865), .I1(1'b1), .CI(n161_2), 
            .O(n158_2), .CO(n159_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i9  (.I0(n867), .I1(n1261), .CI(n168_2), 
            .O(n160_2), .CO(n161_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i8  (.I0(n869), .I1(n1272), .CI(n176_2), 
            .O(n167_2), .CO(n168_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i5  (.I0(n198), .I1(n1277), .CI(n151), 
            .O(n171_2), .CO(n172_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i1  (.I0(\r_mipi_rx_data_1P[30] ), .I1(n1280), 
            .CI(1'b0), .O(n173_2), .CO(n174_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i7  (.I0(n871), .I1(n1282), .CI(n180_2), 
            .O(n175_2), .CO(n176_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i6  (.I0(n873), .I1(n1288), .CI(n199), 
            .O(n179_2), .CO(n180_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i5  (.I0(n875_2), .I1(n1309), .CI(n201), 
            .O(n198), .CO(n199)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i4  (.I0(n877), .I1(n1312), .CI(n203), 
            .O(n200), .CO(n201)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i3  (.I0(n879), .I1(n1315), .CI(n205), 
            .O(n202), .CO(n203)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_70/add_2/i2  (.I0(n881), .I1(n1318), .CI(n416), 
            .O(n204), .CO(n205)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_109/add_2/i11  (.I0(n225), .I1(1'b1), .CI(n208), 
            .O(n206)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_109/add_2/i10  (.I0(n226), .I1(1'b1), .CI(n210), 
            .O(n207), .CO(n208)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_109/add_2/i9  (.I0(n324), .I1(1'b1), .CI(n212), 
            .O(n209), .CO(n210)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_109/add_2/i8  (.I0(n326), .I1(\r_mipi_rx_data_1P[9] ), 
            .CI(n214), .O(n211), .CO(n212)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_109/add_2/i7  (.I0(n330), .I1(\r_mipi_rx_data_1P[8] ), 
            .CI(n216), .O(n213), .CO(n214)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_109/add_2/i6  (.I0(n332), .I1(\r_mipi_rx_data_1P[7] ), 
            .CI(n218), .O(n215), .CO(n216)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_109/add_2/i5  (.I0(n336), .I1(\r_mipi_rx_data_1P[6] ), 
            .CI(n220), .O(n217), .CO(n218)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_109/add_2/i4  (.I0(n338), .I1(\r_mipi_rx_data_1P[5] ), 
            .CI(n222), .O(n219), .CO(n220)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_109/add_2/i3  (.I0(n342), .I1(\r_mipi_rx_data_1P[4] ), 
            .CI(n224), .O(n221), .CO(n222)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_109/add_2/i2  (.I0(n344), .I1(\r_mipi_rx_data_1P[3] ), 
            .CI(n414), .O(n223), .CO(n224)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_109/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_109/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i11  (.I0(n228), .I1(1'b1), .CI(n227), 
            .O(n225)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_106/add_2/i10  (.I0(n229), .I1(1'b1), .CI(n325), 
            .O(n226), .CO(n227)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_55/add_2/i11  (.I0(1'b0), .I1(1'b1), .CI(n230), 
            .O(n228)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_55/add_2/i10  (.I0(\r_mipi_rx_data_1P[9] ), 
            .I1(1'b1), .CI(n232), .O(n229), .CO(n230)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_55/add_2/i9  (.I0(\r_mipi_rx_data_1P[8] ), 
            .I1(1'b1), .CI(n234), .O(n231), .CO(n232)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_55/add_2/i8  (.I0(\r_mipi_rx_data_1P[7] ), 
            .I1(\r_mipi_rx_data_1P[9] ), .CI(n236), .O(n233), .CO(n234)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_55/add_2/i7  (.I0(\r_mipi_rx_data_1P[6] ), 
            .I1(\r_mipi_rx_data_1P[8] ), .CI(n238), .O(n235), .CO(n236)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_55/add_2/i6  (.I0(\r_mipi_rx_data_1P[5] ), 
            .I1(\r_mipi_rx_data_1P[7] ), .CI(n240), .O(n237), .CO(n238)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_55/add_2/i5  (.I0(\r_mipi_rx_data_1P[4] ), 
            .I1(\r_mipi_rx_data_1P[6] ), .CI(n242), .O(n239), .CO(n240)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_55/add_2/i4  (.I0(\r_mipi_rx_data_1P[3] ), 
            .I1(\r_mipi_rx_data_1P[5] ), .CI(n244), .O(n241), .CO(n242)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_55/add_2/i3  (.I0(\r_mipi_rx_data_1P[2] ), 
            .I1(\r_mipi_rx_data_1P[4] ), .CI(n246), .O(n243), .CO(n244)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_55/add_2/i2  (.I0(\r_mipi_rx_data_1P[1] ), 
            .I1(\r_mipi_rx_data_1P[3] ), .CI(n410), .O(n245), .CO(n246)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i11  (.I0(n266), .I1(1'b1), .CI(n249), 
            .O(n247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_49/add_2/i10  (.I0(n267), .I1(1'b1), .CI(n251), 
            .O(n248), .CO(n249)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_49/add_2/i9  (.I0(n269), .I1(1'b1), .CI(n253), 
            .O(n250), .CO(n251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_49/add_2/i8  (.I0(n271_2), .I1(\r_mipi_rx_data_1P[19] ), 
            .CI(n255), .O(n252), .CO(n253)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i7  (.I0(n273), .I1(\r_mipi_rx_data_1P[18] ), 
            .CI(n257), .O(n254), .CO(n255)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i6  (.I0(n275), .I1(\r_mipi_rx_data_1P[17] ), 
            .CI(n259), .O(n256), .CO(n257)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i5  (.I0(n277), .I1(\r_mipi_rx_data_1P[16] ), 
            .CI(n261), .O(n258), .CO(n259)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i4  (.I0(n279), .I1(\r_mipi_rx_data_1P[15] ), 
            .CI(n263), .O(n260), .CO(n261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i3  (.I0(n281), .I1(\r_mipi_rx_data_1P[14] ), 
            .CI(n265), .O(n262), .CO(n263)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i2  (.I0(n283), .I1(\r_mipi_rx_data_1P[13] ), 
            .CI(n408), .O(n264), .CO(n265)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i11  (.I0(n285), .I1(1'b1), .CI(n268), 
            .O(n266)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_46/add_2/i10  (.I0(n286), .I1(1'b1), .CI(n270), 
            .O(n267), .CO(n268)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_46/add_2/i9  (.I0(n288), .I1(\r_mipi_rx_data_1P[19] ), 
            .CI(n272), .O(n269), .CO(n270)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i8  (.I0(n308), .I1(\r_mipi_rx_data_1P[18] ), 
            .CI(n274), .O(n271_2), .CO(n272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i7  (.I0(n322), .I1(\r_mipi_rx_data_1P[17] ), 
            .CI(n276), .O(n273), .CO(n274)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i6  (.I0(n328), .I1(\r_mipi_rx_data_1P[16] ), 
            .CI(n278), .O(n275), .CO(n276)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i5  (.I0(n334), .I1(\r_mipi_rx_data_1P[15] ), 
            .CI(n280), .O(n277), .CO(n278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i4  (.I0(n340), .I1(\r_mipi_rx_data_1P[14] ), 
            .CI(n282), .O(n279), .CO(n280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i3  (.I0(n346), .I1(\r_mipi_rx_data_1P[13] ), 
            .CI(n284), .O(n281), .CO(n282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i2  (.I0(n352), .I1(\r_mipi_rx_data_1P[12] ), 
            .CI(n406), .O(n283), .CO(n284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_43/add_2/i11  (.I0(1'b0), .I1(1'b1), .CI(n287), 
            .O(n285)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_43/add_2/i10  (.I0(\r_mipi_rx_data_1P[19] ), 
            .I1(1'b1), .CI(n289), .O(n286), .CO(n287)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_43/add_2/i9  (.I0(\r_mipi_rx_data_1P[18] ), 
            .I1(1'b1), .CI(n309), .O(n288), .CO(n289)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_43/add_2/i8  (.I0(\r_mipi_rx_data_1P[17] ), 
            .I1(\r_mipi_rx_data_1P[19] ), .CI(n323), .O(n308), .CO(n309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_43/add_2/i7  (.I0(\r_mipi_rx_data_1P[16] ), 
            .I1(\r_mipi_rx_data_1P[18] ), .CI(n329), .O(n322), .CO(n323)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i9  (.I0(n231), .I1(\r_mipi_rx_data_1P[9] ), 
            .CI(n327), .O(n324), .CO(n325)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i8  (.I0(n233), .I1(\r_mipi_rx_data_1P[8] ), 
            .CI(n331), .O(n326), .CO(n327)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_43/add_2/i6  (.I0(\r_mipi_rx_data_1P[15] ), 
            .I1(\r_mipi_rx_data_1P[17] ), .CI(n335), .O(n328), .CO(n329)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i7  (.I0(n235), .I1(\r_mipi_rx_data_1P[7] ), 
            .CI(n333), .O(n330), .CO(n331)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i6  (.I0(n237), .I1(\r_mipi_rx_data_1P[6] ), 
            .CI(n337), .O(n332), .CO(n333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_43/add_2/i5  (.I0(\r_mipi_rx_data_1P[14] ), 
            .I1(\r_mipi_rx_data_1P[16] ), .CI(n341), .O(n334), .CO(n335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i5  (.I0(n239), .I1(\r_mipi_rx_data_1P[5] ), 
            .CI(n339), .O(n336), .CO(n337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i4  (.I0(n241), .I1(\r_mipi_rx_data_1P[4] ), 
            .CI(n343), .O(n338), .CO(n339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_43/add_2/i4  (.I0(\r_mipi_rx_data_1P[13] ), 
            .I1(\r_mipi_rx_data_1P[15] ), .CI(n347), .O(n340), .CO(n341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i3  (.I0(n243), .I1(\r_mipi_rx_data_1P[3] ), 
            .CI(n345), .O(n342), .CO(n343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_106/add_2/i2  (.I0(n245), .I1(\r_mipi_rx_data_1P[2] ), 
            .CI(n412), .O(n344), .CO(n345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(159)
    defparam \inst_line_buf/sub_106/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_106/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_43/add_2/i3  (.I0(\r_mipi_rx_data_1P[12] ), 
            .I1(\r_mipi_rx_data_1P[14] ), .CI(n353), .O(n346), .CO(n347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/add_66/i1  (.I0(n173_2), .I1(n1482), .CI(1'b0), 
            .O(n348), .CO(n349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i1  (.I0(\r_mipi_rx_data_1P[10] ), .I1(n1484), 
            .CI(1'b0), .O(n350), .CO(n351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_43/add_2/i2  (.I0(\r_mipi_rx_data_1P[11] ), 
            .I1(\r_mipi_rx_data_1P[13] ), .CI(n404), .O(n352), .CO(n353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_97/add_2/i11  (.I0(n945_2), .I1(1'b1), .CI(n360), 
            .O(n354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i1  (.I0(n350), .I1(n1490), .CI(1'b0), 
            .O(n355), .CO(n356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_19/add_2/i1  (.I0(\r_mipi_rx_data_1P[30] ), 
            .I1(\r_mipi_rx_data_1P[32] ), .CI(n2425), .O(n357), .CO(n358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_97/add_2/i10  (.I0(n946), .I1(1'b1), .CI(n362), 
            .O(n359), .CO(n360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_97/add_2/i9  (.I0(n948), .I1(1'b1), .CI(n366_2), 
            .O(n361), .CO(n362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_25/add_2/i1  (.I0(n369_2), .I1(\r_mipi_rx_data_1P[32] ), 
            .CI(n2426), .O(n363), .CO(n364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_97/add_2/i8  (.I0(n950_2), .I1(n1498), .CI(n368_2), 
            .O(n365_2), .CO(n366_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_97/add_2/i7  (.I0(n952), .I1(n1501), .CI(n372_2), 
            .O(n367_2), .CO(n368_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_22/add_2/i1  (.I0(n357), .I1(\r_mipi_rx_data_1P[31] ), 
            .CI(n2427), .O(n369_2), .CO(n370_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_97/add_2/i6  (.I0(n954), .I1(n1506), .CI(n395), 
            .O(n371_2), .CO(n372_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_31/add_2/i1  (.I0(\r_mipi_rx_data_1P[20] ), 
            .I1(\r_mipi_rx_data_1P[22] ), .CI(n2428), .O(n373_2), .CO(n374_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_97/add_2/i5  (.I0(n956), .I1(n1533), .CI(n940_2), 
            .O(n394), .CO(n395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_37/add_2/i1  (.I0(n419), .I1(\r_mipi_rx_data_1P[22] ), 
            .CI(n2429), .O(n401), .CO(n402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_37/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_37/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_43/add_2/i1  (.I0(\r_mipi_rx_data_1P[10] ), 
            .I1(\r_mipi_rx_data_1P[12] ), .CI(n2430), .O(n403), .CO(n404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_43/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_43/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_46/add_2/i1  (.I0(n403), .I1(\r_mipi_rx_data_1P[11] ), 
            .CI(n2431), .O(n405), .CO(n406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_46/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_46/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_49/add_2/i1  (.I0(n405), .I1(\r_mipi_rx_data_1P[12] ), 
            .CI(n2432), .O(n407), .CO(n408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(144)
    defparam \inst_line_buf/sub_49/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_49/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_55/add_2/i1  (.I0(\r_mipi_rx_data_1P[0] ), 
            .I1(\r_mipi_rx_data_1P[2] ), .CI(n2433), .O(n409), .CO(n410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_55/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_55/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_58/add_2/i1  (.I0(n409), .I1(\r_mipi_rx_data_1P[1] ), 
            .CI(n2434), .O(n411), .CO(n412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_58/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_58/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_61/add_2/i1  (.I0(n411), .I1(\r_mipi_rx_data_1P[2] ), 
            .CI(n2435), .O(n413), .CO(n414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(147)
    defparam \inst_line_buf/sub_61/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_61/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_70/add_2/i1  (.I0(n357), .I1(n1548), .CI(n2436), 
            .O(n415), .CO(n416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_70/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_70/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i1  (.I0(n415), .I1(n1550), .CI(n2437), 
            .O(n417), .CO(n418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_82/add_2/i1  (.I0(n373_2), .I1(\r_mipi_rx_data_1P[21] ), 
            .CI(n2438), .O(n419), .CO(n420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i1 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_94/add_2/i1  (.I0(n403), .I1(n1553), .CI(n2439), 
            .O(n421), .CO(n422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_97/add_2/i1  (.I0(n421), .I1(n1555), .CI(n2440), 
            .O(n423), .CO(n424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i1 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i1 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_34/add_2/i2  (.I0(n824), .I1(\r_mipi_rx_data_1P[22] ), 
            .CI(n420), .O(n805), .CO(n806)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_34/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_34/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_31/add_2/i11  (.I0(1'b0), .I1(1'b1), .CI(n809), 
            .O(n807)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_31/add_2/i10  (.I0(\r_mipi_rx_data_1P[29] ), 
            .I1(1'b1), .CI(n811), .O(n808), .CO(n809)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_31/add_2/i9  (.I0(\r_mipi_rx_data_1P[28] ), 
            .I1(1'b1), .CI(n813), .O(n810), .CO(n811)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_31/add_2/i8  (.I0(\r_mipi_rx_data_1P[27] ), 
            .I1(\r_mipi_rx_data_1P[29] ), .CI(n815), .O(n812), .CO(n813)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_31/add_2/i7  (.I0(\r_mipi_rx_data_1P[26] ), 
            .I1(\r_mipi_rx_data_1P[28] ), .CI(n817), .O(n814), .CO(n815)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_31/add_2/i6  (.I0(\r_mipi_rx_data_1P[25] ), 
            .I1(\r_mipi_rx_data_1P[27] ), .CI(n819), .O(n816), .CO(n817)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_31/add_2/i5  (.I0(\r_mipi_rx_data_1P[24] ), 
            .I1(\r_mipi_rx_data_1P[26] ), .CI(n821), .O(n818), .CO(n819)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_31/add_2/i4  (.I0(\r_mipi_rx_data_1P[23] ), 
            .I1(\r_mipi_rx_data_1P[25] ), .CI(n823), .O(n820), .CO(n821)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_31/add_2/i3  (.I0(\r_mipi_rx_data_1P[22] ), 
            .I1(\r_mipi_rx_data_1P[24] ), .CI(n825), .O(n822), .CO(n823)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_31/add_2/i2  (.I0(\r_mipi_rx_data_1P[21] ), 
            .I1(\r_mipi_rx_data_1P[23] ), .CI(n374_2), .O(n824), .CO(n825)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(141)
    defparam \inst_line_buf/sub_31/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_31/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i11  (.I0(n864), .I1(1'b1), .CI(n828), 
            .O(n826)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_22/add_2/i10  (.I0(n865), .I1(1'b1), .CI(n830), 
            .O(n827), .CO(n828)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_22/add_2/i9  (.I0(n867), .I1(\r_mipi_rx_data_1P[39] ), 
            .CI(n832), .O(n829), .CO(n830)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i8  (.I0(n869), .I1(\r_mipi_rx_data_1P[38] ), 
            .CI(n834), .O(n831), .CO(n832)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i7  (.I0(n871), .I1(\r_mipi_rx_data_1P[37] ), 
            .CI(n836), .O(n833), .CO(n834)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i6  (.I0(n873), .I1(\r_mipi_rx_data_1P[36] ), 
            .CI(n838), .O(n835), .CO(n836)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i5  (.I0(n875_2), .I1(\r_mipi_rx_data_1P[35] ), 
            .CI(n840), .O(n837), .CO(n838)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i4  (.I0(n877), .I1(\r_mipi_rx_data_1P[34] ), 
            .CI(n842), .O(n839), .CO(n840)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i3  (.I0(n879), .I1(\r_mipi_rx_data_1P[33] ), 
            .CI(n844), .O(n841), .CO(n842)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_22/add_2/i2  (.I0(n881), .I1(\r_mipi_rx_data_1P[32] ), 
            .CI(n370_2), .O(n843), .CO(n844)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_22/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_22/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_25/add_2/i11  (.I0(n826), .I1(1'b1), .CI(n847), 
            .O(n845)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_25/add_2/i10  (.I0(n827), .I1(1'b1), .CI(n849), 
            .O(n846), .CO(n847)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_25/add_2/i9  (.I0(n829), .I1(1'b1), .CI(n851), 
            .O(n848), .CO(n849)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_25/add_2/i8  (.I0(n831), .I1(\r_mipi_rx_data_1P[39] ), 
            .CI(n853), .O(n850), .CO(n851)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_25/add_2/i7  (.I0(n833), .I1(\r_mipi_rx_data_1P[38] ), 
            .CI(n855), .O(n852), .CO(n853)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_25/add_2/i6  (.I0(n835), .I1(\r_mipi_rx_data_1P[37] ), 
            .CI(n857), .O(n854), .CO(n855)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_25/add_2/i5  (.I0(n837), .I1(\r_mipi_rx_data_1P[36] ), 
            .CI(n859), .O(n856), .CO(n857)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_25/add_2/i4  (.I0(n839), .I1(\r_mipi_rx_data_1P[35] ), 
            .CI(n861), .O(n858), .CO(n859)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_25/add_2/i3  (.I0(n841), .I1(\r_mipi_rx_data_1P[34] ), 
            .CI(n863), .O(n860), .CO(n861)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_25/add_2/i2  (.I0(n843), .I1(\r_mipi_rx_data_1P[33] ), 
            .CI(n364), .O(n862), .CO(n863)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_25/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_25/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_19/add_2/i11  (.I0(1'b0), .I1(1'b1), .CI(n866), 
            .O(n864)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_19/add_2/i10  (.I0(\r_mipi_rx_data_1P[39] ), 
            .I1(1'b1), .CI(n868), .O(n865), .CO(n866)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_19/add_2/i9  (.I0(\r_mipi_rx_data_1P[38] ), 
            .I1(1'b1), .CI(n870), .O(n867), .CO(n868)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_19/add_2/i8  (.I0(\r_mipi_rx_data_1P[37] ), 
            .I1(\r_mipi_rx_data_1P[39] ), .CI(n872), .O(n869), .CO(n870)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_19/add_2/i7  (.I0(\r_mipi_rx_data_1P[36] ), 
            .I1(\r_mipi_rx_data_1P[38] ), .CI(n874_2), .O(n871), .CO(n872)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_19/add_2/i6  (.I0(\r_mipi_rx_data_1P[35] ), 
            .I1(\r_mipi_rx_data_1P[37] ), .CI(n876), .O(n873), .CO(n874_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_19/add_2/i5  (.I0(\r_mipi_rx_data_1P[34] ), 
            .I1(\r_mipi_rx_data_1P[36] ), .CI(n878), .O(n875_2), .CO(n876)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_19/add_2/i4  (.I0(\r_mipi_rx_data_1P[33] ), 
            .I1(\r_mipi_rx_data_1P[35] ), .CI(n880), .O(n877), .CO(n878)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_19/add_2/i3  (.I0(\r_mipi_rx_data_1P[32] ), 
            .I1(\r_mipi_rx_data_1P[34] ), .CI(n882), .O(n879), .CO(n880)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_19/add_2/i2  (.I0(\r_mipi_rx_data_1P[31] ), 
            .I1(\r_mipi_rx_data_1P[33] ), .CI(n358), .O(n881), .CO(n882)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(138)
    defparam \inst_line_buf/sub_19/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_19/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/add_90/i11  (.I0(n903), .I1(1'b0), .CI(n885_2), 
            .O(n883)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i10  (.I0(n902), .I1(1'b0), .CI(n887), 
            .O(n884), .CO(n885_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i9  (.I0(n904), .I1(1'b0), .CI(n889), 
            .O(n886), .CO(n887)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i8  (.I0(n906), .I1(n2071), .CI(n891), 
            .O(n888), .CO(n889)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i7  (.I0(n908), .I1(n2074), .CI(n893), 
            .O(n890_2), .CO(n891)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i6  (.I0(n910_2), .I1(n2077), .CI(n895_2), 
            .O(n892), .CO(n893)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i5  (.I0(n912), .I1(n2080), .CI(n897), 
            .O(n894), .CO(n895_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i4  (.I0(n914), .I1(n2083), .CI(n899), 
            .O(n896), .CO(n897)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i3  (.I0(n916), .I1(n2086), .CI(n901), 
            .O(n898), .CO(n899)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_90/i2  (.I0(n918), .I1(n2089), .CI(n356), 
            .O(n900_2), .CO(n901)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_90/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_90/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i10  (.I0(\r_mipi_rx_data_1P[19] ), .I1(1'b0), 
            .CI(n905_2), .O(n902), .CO(n2441)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i9  (.I0(\r_mipi_rx_data_1P[18] ), .I1(n2092), 
            .CI(n907), .O(n904), .CO(n905_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i8  (.I0(\r_mipi_rx_data_1P[17] ), .I1(n2094), 
            .CI(n909), .O(n906), .CO(n907)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i7  (.I0(\r_mipi_rx_data_1P[16] ), .I1(n2096), 
            .CI(n911), .O(n908), .CO(n909)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i6  (.I0(\r_mipi_rx_data_1P[15] ), .I1(n2098), 
            .CI(n913), .O(n910_2), .CO(n911)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i5  (.I0(\r_mipi_rx_data_1P[14] ), .I1(n2100), 
            .CI(n915_2), .O(n912), .CO(n913)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i4  (.I0(\r_mipi_rx_data_1P[13] ), .I1(n2102), 
            .CI(n917), .O(n914), .CO(n915_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i3  (.I0(\r_mipi_rx_data_1P[12] ), .I1(n2104), 
            .CI(n919), .O(n916), .CO(n917)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_88/i2  (.I0(\r_mipi_rx_data_1P[11] ), .I1(n2106), 
            .CI(n351), .O(n918), .CO(n919)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(155)
    defparam \inst_line_buf/add_88/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_88/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i11  (.I0(n961), .I1(1'b0), .CI(n922), 
            .O(n920_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i10  (.I0(n960), .I1(1'b0), .CI(n924), 
            .O(n921), .CO(n922)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i9  (.I0(n962), .I1(1'b0), .CI(n926), 
            .O(n923), .CO(n924)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i8  (.I0(n964), .I1(n2115), .CI(n928), 
            .O(n925_2), .CO(n926)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i7  (.I0(n966), .I1(n2118), .CI(n930_2), 
            .O(n927), .CO(n928)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i6  (.I0(n968), .I1(n2121), .CI(n932), 
            .O(n929), .CO(n930_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i5  (.I0(n970), .I1(n2124), .CI(n934), 
            .O(n931), .CO(n932)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i4  (.I0(n972), .I1(n2127), .CI(n936), 
            .O(n933), .CO(n934)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i3  (.I0(n974), .I1(n2130), .CI(n938), 
            .O(n935_2), .CO(n936)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_66/i2  (.I0(n976), .I1(n2133), .CI(n349), 
            .O(n937), .CO(n938)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_66/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_66/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_97/add_2/i4  (.I0(n958), .I1(n2136), .CI(n942), 
            .O(n939), .CO(n940_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_97/add_2/i3  (.I0(n1030), .I1(n2139), .CI(n944), 
            .O(n941), .CO(n942)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_97/add_2/i2  (.I0(n1032), .I1(n2142), .CI(n424), 
            .O(n943), .CO(n944)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_97/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_97/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i11  (.I0(n285), .I1(1'b1), .CI(n947), 
            .O(n945_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i10  (.I0(n286), .I1(1'b1), .CI(n949), 
            .O(n946), .CO(n947)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i9  (.I0(n288), .I1(n2146), .CI(n951), 
            .O(n948), .CO(n949)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i8  (.I0(n308), .I1(n2148), .CI(n953), 
            .O(n950_2), .CO(n951)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i7  (.I0(n322), .I1(n2150), .CI(n955_2), 
            .O(n952), .CO(n953)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i6  (.I0(n328), .I1(n2152), .CI(n957), 
            .O(n954), .CO(n955_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i5  (.I0(n334), .I1(n2154), .CI(n959), 
            .O(n956), .CO(n957)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i4  (.I0(n340), .I1(n2156), .CI(n1031), 
            .O(n958), .CO(n959)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i10  (.I0(\r_mipi_rx_data_1P[39] ), .I1(1'b0), 
            .CI(n963), .O(n960), .CO(n2442)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i9  (.I0(\r_mipi_rx_data_1P[38] ), .I1(n2159), 
            .CI(n965), .O(n962), .CO(n963)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i8  (.I0(\r_mipi_rx_data_1P[37] ), .I1(n2161), 
            .CI(n967), .O(n964), .CO(n965)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i7  (.I0(\r_mipi_rx_data_1P[36] ), .I1(n2163), 
            .CI(n969), .O(n966), .CO(n967)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i6  (.I0(\r_mipi_rx_data_1P[35] ), .I1(n2165), 
            .CI(n971), .O(n968), .CO(n969)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i5  (.I0(\r_mipi_rx_data_1P[34] ), .I1(n2167), 
            .CI(n973), .O(n970), .CO(n971)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i4  (.I0(\r_mipi_rx_data_1P[33] ), .I1(n2169), 
            .CI(n975), .O(n972), .CO(n973)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i3  (.I0(\r_mipi_rx_data_1P[32] ), .I1(n2171), 
            .CI(n977), .O(n974), .CO(n975)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/add_64/i2  (.I0(\r_mipi_rx_data_1P[31] ), .I1(n2173), 
            .CI(n174_2), .O(n976), .CO(n977)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(149)
    defparam \inst_line_buf/add_64/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/add_64/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i13  (.I0(\r_waddr_1P[12]_2 ), .I1(1'b0), .CI(n980), 
            .O(n978)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i13 .I0_POLARITY = 1'b1;
    defparam \add_81/i13 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i12  (.I0(\r_waddr_1P[11]_2 ), .I1(1'b0), .CI(n996), 
            .O(n979), .CO(n980)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i12 .I0_POLARITY = 1'b1;
    defparam \add_81/i12 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i11  (.I0(\r_waddr_1P[10]_2 ), .I1(1'b0), .CI(n999), 
            .O(n995), .CO(n996)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i11 .I0_POLARITY = 1'b1;
    defparam \add_81/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i10  (.I0(\r_waddr_1P[9]_2 ), .I1(1'b0), .CI(n1001), 
            .O(n998), .CO(n999)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i10 .I0_POLARITY = 1'b1;
    defparam \add_81/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i9  (.I0(\r_waddr_1P[8]_2 ), .I1(1'b0), .CI(n1027), 
            .O(n1000), .CO(n1001)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i9 .I0_POLARITY = 1'b1;
    defparam \add_81/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i8  (.I0(\r_waddr_1P[7]_2 ), .I1(1'b0), .CI(n1029), 
            .O(n1026), .CO(n1027)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i8 .I0_POLARITY = 1'b1;
    defparam \add_81/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i7  (.I0(\r_waddr_1P[6]_2 ), .I1(1'b0), .CI(n1057), 
            .O(n1028), .CO(n1029)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i7 .I0_POLARITY = 1'b1;
    defparam \add_81/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i3  (.I0(n346), .I1(n2221), .CI(n1033), 
            .O(n1030), .CO(n1031)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_94/add_2/i2  (.I0(n352), .I1(n2223), .CI(n422), 
            .O(n1032), .CO(n1033)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(156)
    defparam \inst_line_buf/sub_94/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_94/add_2/i2 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_85/add_2/i11  (.I0(n1053), .I1(1'b1), .CI(n1036), 
            .O(n1034)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_85/add_2/i10  (.I0(n1054), .I1(1'b1), .CI(n1038), 
            .O(n1035), .CO(n1036)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_85/add_2/i9  (.I0(n1065_2), .I1(1'b1), .CI(n1040), 
            .O(n1037), .CO(n1038)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_85/add_2/i8  (.I0(n1067), .I1(\r_mipi_rx_data_1P[29] ), 
            .CI(n1042), .O(n1039), .CO(n1040)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_85/add_2/i7  (.I0(n1071), .I1(\r_mipi_rx_data_1P[28] ), 
            .CI(n1044), .O(n1041), .CO(n1042)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_85/add_2/i6  (.I0(n1073), .I1(\r_mipi_rx_data_1P[27] ), 
            .CI(n1046), .O(n1043), .CO(n1044)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_85/add_2/i5  (.I0(n1075_2), .I1(\r_mipi_rx_data_1P[26] ), 
            .CI(n1048), .O(n1045), .CO(n1046)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_85/add_2/i4  (.I0(n1077), .I1(\r_mipi_rx_data_1P[25] ), 
            .CI(n1050), .O(n1047), .CO(n1048)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_85/add_2/i3  (.I0(n1079), .I1(\r_mipi_rx_data_1P[24] ), 
            .CI(n1052), .O(n1049), .CO(n1050)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_85/add_2/i2  (.I0(n805), .I1(\r_mipi_rx_data_1P[23] ), 
            .CI(n402), .O(n1051), .CO(n1052)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_85/add_2/i2 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_85/add_2/i2 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_82/add_2/i11  (.I0(n807), .I1(1'b1), .CI(n1055), 
            .O(n1053)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_82/add_2/i10  (.I0(n808), .I1(1'b1), .CI(n1066), 
            .O(n1054), .CO(n1055)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i6  (.I0(\r_waddr_1P[5]_2 ), .I1(1'b0), .CI(n1059), 
            .O(n1056), .CO(n1057)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i6 .I0_POLARITY = 1'b1;
    defparam \add_81/i6 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i5  (.I0(\r_waddr_1P[4]_2 ), .I1(1'b0), .CI(n1061), 
            .O(n1058), .CO(n1059)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i5 .I0_POLARITY = 1'b1;
    defparam \add_81/i5 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i4  (.I0(\r_waddr_1P[3]_2 ), .I1(1'b0), .CI(n1063), 
            .O(n1060_2), .CO(n1061)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i4 .I0_POLARITY = 1'b1;
    defparam \add_81/i4 .I1_POLARITY = 1'b1;
    EFX_ADD \add_81/i3  (.I0(\r_waddr_1P[2]_2 ), .I1(1'b0), .CI(n142), 
            .O(n1062), .CO(n1063)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\mipi_pi_top.v(244)
    defparam \add_81/i3 .I0_POLARITY = 1'b1;
    defparam \add_81/i3 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_82/add_2/i9  (.I0(n810), .I1(\r_mipi_rx_data_1P[29] ), 
            .CI(n1068), .O(n1065_2), .CO(n1066)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i9 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_82/add_2/i8  (.I0(n812), .I1(\r_mipi_rx_data_1P[28] ), 
            .CI(n1072), .O(n1067), .CO(n1068)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i8 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_82/add_2/i7  (.I0(n814), .I1(\r_mipi_rx_data_1P[27] ), 
            .CI(n1074), .O(n1071), .CO(n1072)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i7 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_82/add_2/i6  (.I0(n816), .I1(\r_mipi_rx_data_1P[26] ), 
            .CI(n1076), .O(n1073), .CO(n1074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i6 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_82/add_2/i5  (.I0(n818), .I1(\r_mipi_rx_data_1P[25] ), 
            .CI(n1078), .O(n1075_2), .CO(n1076)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i5 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i5 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_82/add_2/i4  (.I0(n820), .I1(\r_mipi_rx_data_1P[24] ), 
            .CI(n1080_2), .O(n1077), .CO(n1078)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i4 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i4 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_82/add_2/i3  (.I0(n822), .I1(\r_mipi_rx_data_1P[23] ), 
            .CI(n806), .O(n1079), .CO(n1080_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(153)
    defparam \inst_line_buf/sub_82/add_2/i3 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_82/add_2/i3 .I1_POLARITY = 1'b0;
    EFX_ADD \inst_line_buf/sub_73/add_2/i11  (.I0(n157), .I1(1'b1), .CI(n1083), 
            .O(n1081)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i11 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i11 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i10  (.I0(n158_2), .I1(1'b1), .CI(n1085_2), 
            .O(n1082), .CO(n1083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i10 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i10 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i9  (.I0(n160_2), .I1(1'b1), .CI(n1087), 
            .O(n1084), .CO(n1085_2)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i9 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i9 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i8  (.I0(n167_2), .I1(n2278), .CI(n1089), 
            .O(n1086), .CO(n1087)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i8 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i8 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i7  (.I0(n175_2), .I1(n2281), .CI(n1091), 
            .O(n1088), .CO(n1089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i7 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i7 .I1_POLARITY = 1'b1;
    EFX_ADD \inst_line_buf/sub_73/add_2/i6  (.I0(n179_2), .I1(n2284), .CI(n172_2), 
            .O(n1090_2), .CO(n1091)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_ADD, I0_POLARITY=1'b1, I1_POLARITY=1'b1 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\line_buf_4_to_6.v(150)
    defparam \inst_line_buf/sub_73/add_2/i6 .I0_POLARITY = 1'b1;
    defparam \inst_line_buf/sub_73/add_2/i6 .I1_POLARITY = 1'b1;
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$2  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[1]_2 , \inst_line_buf/r_mipi_rx_data_1P[0]_2 }), 
            .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , \inst_line_buf/r_mipi_rx_x_2P[9]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[8]_2 , \inst_line_buf/r_mipi_rx_x_2P[7]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[6]_2 , \inst_line_buf/r_mipi_rx_x_2P[5]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[4]_2 , \inst_line_buf/r_mipi_rx_x_2P[3]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[2]_2 , \inst_line_buf/r_mipi_rx_x_2P[1]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[9]_2 , \inst_line_buf/r_mipi_tx_x_1P[8]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[7]_2 , \inst_line_buf/r_mipi_tx_x_1P[6]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[5]_2 , \inst_line_buf/r_mipi_tx_x_1P[4]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[3]_2 , \inst_line_buf/r_mipi_tx_x_1P[2]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[1]_2 , \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), 
            .RDATA({\inst_line_buf/w_mipi_tx_data_3P[1] , \inst_line_buf/w_mipi_tx_data_3P[0] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$2 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[3]_2 , \inst_line_buf/r_mipi_rx_data_1P[2]_2 }), 
            .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , \inst_line_buf/r_mipi_rx_x_2P[9]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[8]_2 , \inst_line_buf/r_mipi_rx_x_2P[7]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[6]_2 , \inst_line_buf/r_mipi_rx_x_2P[5]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[4]_2 , \inst_line_buf/r_mipi_rx_x_2P[3]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[2]_2 , \inst_line_buf/r_mipi_rx_x_2P[1]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[9]_2 , \inst_line_buf/r_mipi_tx_x_1P[8]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[7]_2 , \inst_line_buf/r_mipi_tx_x_1P[6]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[5]_2 , \inst_line_buf/r_mipi_tx_x_1P[4]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[3]_2 , \inst_line_buf/r_mipi_tx_x_1P[2]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[1]_2 , \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), 
            .RDATA({\inst_line_buf/w_mipi_tx_data_3P[3] , \inst_line_buf/w_mipi_tx_data_3P[2] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_dly/ram__D$3  (.WCLK(\mipi_pclk~O ), .RCLK(\mipi_pclk~O ), 
            .WCLKE(1'b1), .WE(\r_waddr_1P[12]_2 ), .RE(n1502), .WDATA({rx_status}), 
            .WADDR({\r_waddr_1P[11]_2 , \r_waddr_1P[10]_2 , \r_waddr_1P[9]_2 , 
            \r_waddr_1P[8]_2 , \r_waddr_1P[7]_2 , \r_waddr_1P[6]_2 , \r_waddr_1P[5]_2 , 
            \r_waddr_1P[4]_2 , \r_waddr_1P[3]_2 , \r_waddr_1P[2]_2 , \r_waddr_1P[1]_2 , 
            \r_waddr_1P[0]_2 }), .RADDR({\r_raddr_1P[11]_2 , \r_raddr_1P[10]_2 , 
            \r_raddr_1P[9]_2 , \r_raddr_1P[8]_2 , \r_raddr_1P[7]_2 , \r_raddr_1P[6]_2 , 
            \r_raddr_1P[5]_2 , \r_raddr_1P[4]_2 , \r_raddr_1P[3]_2 , \r_raddr_1P[2]_2 , 
            \r_raddr_1P[1]_2 , \r_raddr_1P[0]_2 }), .RDATA({\inst_dly/n28 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_dly/ram__D$3 .READ_WIDTH = 1;
    defparam \inst_dly/ram__D$3 .WRITE_WIDTH = 1;
    defparam \inst_dly/ram__D$3 .WCLK_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$3 .WCLKE_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$3 .WE_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$3 .RCLK_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$3 .RE_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$3 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$3 .OUTPUT_REG = 1'b0;
    defparam \inst_dly/ram__D$3 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[5]_2 , \inst_line_buf/r_mipi_rx_data_1P[4]_2 }), 
            .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , \inst_line_buf/r_mipi_rx_x_2P[9]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[8]_2 , \inst_line_buf/r_mipi_rx_x_2P[7]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[6]_2 , \inst_line_buf/r_mipi_rx_x_2P[5]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[4]_2 , \inst_line_buf/r_mipi_rx_x_2P[3]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[2]_2 , \inst_line_buf/r_mipi_rx_x_2P[1]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[9]_2 , \inst_line_buf/r_mipi_tx_x_1P[8]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[7]_2 , \inst_line_buf/r_mipi_tx_x_1P[6]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[5]_2 , \inst_line_buf/r_mipi_tx_x_1P[4]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[3]_2 , \inst_line_buf/r_mipi_tx_x_1P[2]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[1]_2 , \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), 
            .RDATA({\inst_line_buf/w_mipi_tx_data_3P[5] , \inst_line_buf/w_mipi_tx_data_3P[4] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$b12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[7]_2 , \inst_line_buf/r_mipi_rx_data_1P[6]_2 }), 
            .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , \inst_line_buf/r_mipi_rx_x_2P[9]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[8]_2 , \inst_line_buf/r_mipi_rx_x_2P[7]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[6]_2 , \inst_line_buf/r_mipi_rx_x_2P[5]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[4]_2 , \inst_line_buf/r_mipi_rx_x_2P[3]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[2]_2 , \inst_line_buf/r_mipi_rx_x_2P[1]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[9]_2 , \inst_line_buf/r_mipi_tx_x_1P[8]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[7]_2 , \inst_line_buf/r_mipi_tx_x_1P[6]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[5]_2 , \inst_line_buf/r_mipi_tx_x_1P[4]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[3]_2 , \inst_line_buf/r_mipi_tx_x_1P[2]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[1]_2 , \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), 
            .RDATA({\inst_line_buf/w_mipi_tx_data_3P[7] , \inst_line_buf/w_mipi_tx_data_3P[6] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$c12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[9]_2 , \inst_line_buf/r_mipi_rx_data_1P[8]_2 }), 
            .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , \inst_line_buf/r_mipi_rx_x_2P[9]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[8]_2 , \inst_line_buf/r_mipi_rx_x_2P[7]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[6]_2 , \inst_line_buf/r_mipi_rx_x_2P[5]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[4]_2 , \inst_line_buf/r_mipi_rx_x_2P[3]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[2]_2 , \inst_line_buf/r_mipi_rx_x_2P[1]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[9]_2 , \inst_line_buf/r_mipi_tx_x_1P[8]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[7]_2 , \inst_line_buf/r_mipi_tx_x_1P[6]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[5]_2 , \inst_line_buf/r_mipi_tx_x_1P[4]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[3]_2 , \inst_line_buf/r_mipi_tx_x_1P[2]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[1]_2 , \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), 
            .RDATA({\inst_line_buf/w_mipi_tx_data_3P[9] , \inst_line_buf/w_mipi_tx_data_3P[8] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$d12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[11]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[10]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[11] , 
            \inst_line_buf/w_mipi_tx_data_3P[10] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$e12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[13]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[12]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[13] , 
            \inst_line_buf/w_mipi_tx_data_3P[12] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$f12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[15]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[14]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[15] , 
            \inst_line_buf/w_mipi_tx_data_3P[14] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$g12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[17]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[16]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[17] , 
            \inst_line_buf/w_mipi_tx_data_3P[16] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$h12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[19]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[18]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[19] , 
            \inst_line_buf/w_mipi_tx_data_3P[18] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$i12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[21]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[20]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[21] , 
            \inst_line_buf/w_mipi_tx_data_3P[20] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$j12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[23]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[22]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[23] , 
            \inst_line_buf/w_mipi_tx_data_3P[22] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$k12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[25]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[24]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[25] , 
            \inst_line_buf/w_mipi_tx_data_3P[24] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$l12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[27]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[26]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[27] , 
            \inst_line_buf/w_mipi_tx_data_3P[26] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$m12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[29]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[28]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[29] , 
            \inst_line_buf/w_mipi_tx_data_3P[28] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$n12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[31]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[30]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[31] , 
            \inst_line_buf/w_mipi_tx_data_3P[30] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$o12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[33]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[32]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[33] , 
            \inst_line_buf/w_mipi_tx_data_3P[32] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$p12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[35]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[34]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[35] , 
            \inst_line_buf/w_mipi_tx_data_3P[34] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$q12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[37]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[36]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[37] , 
            \inst_line_buf/w_mipi_tx_data_3P[36] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$r12 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1  (.WCLK(\mipi_pclk~O ), 
            .RCLK(\mipi_pclk~O ), .WCLKE(1'b1), .WE(\inst_line_buf/r_mipi_rx_valid_1P_2 ), 
            .RE(1'b1), .WDATA({\inst_line_buf/r_mipi_rx_data_1P[39]_2 , 
            \inst_line_buf/r_mipi_rx_data_1P[38]_2 }), .WADDR({\inst_line_buf/r_mipi_rx_x_2P[10]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[9]_2 , \inst_line_buf/r_mipi_rx_x_2P[8]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[7]_2 , \inst_line_buf/r_mipi_rx_x_2P[6]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[5]_2 , \inst_line_buf/r_mipi_rx_x_2P[4]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[3]_2 , \inst_line_buf/r_mipi_rx_x_2P[2]_2 , 
            \inst_line_buf/r_mipi_rx_x_2P[1]_2 , \inst_line_buf/r_mipi_rx_x_2P[0]_2 }), 
            .RADDR({\inst_line_buf/r_mipi_tx_x_1P[10]_2 , \inst_line_buf/r_mipi_tx_x_1P[9]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[8]_2 , \inst_line_buf/r_mipi_tx_x_1P[7]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[6]_2 , \inst_line_buf/r_mipi_tx_x_1P[5]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[4]_2 , \inst_line_buf/r_mipi_tx_x_1P[3]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[2]_2 , \inst_line_buf/r_mipi_tx_x_1P[1]_2 , 
            \inst_line_buf/r_mipi_tx_x_1P[0]_2 }), .RDATA({\inst_line_buf/w_mipi_tx_data_3P[39] , 
            \inst_line_buf/w_mipi_tx_data_3P[38] })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=2, WRITE_WIDTH=2, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b1, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b1, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .READ_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .WRITE_WIDTH = 2;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .WCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .WCLKE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .WE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .RCLK_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .RE_POLARITY = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .OUTPUT_REG = 1'b1;
    defparam \inst_line_buf/inst_simple_dual_port_ram/ram__D$s1 .WRITE_MODE = "READ_FIRST";
    EFX_RAM_5K \inst_dly/ram__D$0  (.WCLK(\mipi_pclk~O ), .RCLK(\mipi_pclk~O ), 
            .WCLKE(1'b1), .WE(\r_waddr_1P[12]_2 ), .RE(n1504), .WDATA({rx_status}), 
            .WADDR({\r_waddr_1P[11]_2 , \r_waddr_1P[10]_2 , \r_waddr_1P[9]_2 , 
            \r_waddr_1P[8]_2 , \r_waddr_1P[7]_2 , \r_waddr_1P[6]_2 , \r_waddr_1P[5]_2 , 
            \r_waddr_1P[4]_2 , \r_waddr_1P[3]_2 , \r_waddr_1P[2]_2 , \r_waddr_1P[1]_2 , 
            \r_waddr_1P[0]_2 }), .RADDR({\r_raddr_1P[11]_2 , \r_raddr_1P[10]_2 , 
            \r_raddr_1P[9]_2 , \r_raddr_1P[8]_2 , \r_raddr_1P[7]_2 , \r_raddr_1P[6]_2 , 
            \r_raddr_1P[5]_2 , \r_raddr_1P[4]_2 , \r_raddr_1P[3]_2 , \r_raddr_1P[2]_2 , 
            \r_raddr_1P[1]_2 , \r_raddr_1P[0]_2 }), .RDATA({\inst_dly/n29 })) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_RAM_5K, READ_WIDTH=1, WRITE_WIDTH=1, WCLK_POLARITY=1'b1, WCLKE_POLARITY=1'b1, WE_POLARITY=1'b0, RCLK_POLARITY=1'b1, RE_POLARITY=1'b1, OUTPUT_REG=1'b0, WRITE_MODE="READ_FIRST", INIT_0=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_1=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_2=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_3=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_4=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_5=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_6=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_7=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_8=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_9=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_A=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_B=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_C=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_D=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_E=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_F=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_10=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_11=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_12=256'h0000000000000000000000000000000000000000000000000000000000000000, INIT_13=256'h0000000000000000000000000000000000000000000000000000000000000000, PRESERVE_USER_INIT=1'b0 */ ;   // C:/Users\sanas\OneDrive\Documents\t120_bridge\bridge_T120\simple_dual_port_ram.v(31)
    defparam \inst_dly/ram__D$0 .READ_WIDTH = 1;
    defparam \inst_dly/ram__D$0 .WRITE_WIDTH = 1;
    defparam \inst_dly/ram__D$0 .WCLK_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$0 .WCLKE_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$0 .WE_POLARITY = 1'b0;
    defparam \inst_dly/ram__D$0 .RCLK_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$0 .RE_POLARITY = 1'b1;
    defparam \inst_dly/ram__D$0 .INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    defparam \inst_dly/ram__D$0 .OUTPUT_REG = 1'b0;
    defparam \inst_dly/ram__D$0 .WRITE_MODE = "READ_FIRST";
    EFX_LUT4 LUT__3517 (.I0(\key1_counter[8] ), .I1(\key1_counter[9] ), 
            .I2(\key1_counter[14] ), .I3(\key1_counter[15] ), .O(n2332)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3517.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3518 (.I0(\key1_counter[10] ), .I1(\key1_counter[11] ), 
            .I2(\key1_counter[12] ), .I3(\key1_counter[13] ), .O(n2333)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3518.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3519 (.I0(n2333), .I1(\key1_counter[15] ), .I2(\key1_counter[14] ), 
            .I3(key1), .O(n2334)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h00bf */ ;
    defparam LUT__3519.LUTMASK = 16'h00bf;
    EFX_LUT4 LUT__3520 (.I0(\key1_counter[7] ), .I1(n2331), .I2(n2332), 
            .I3(n2334), .O(n271)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__3520.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__3521 (.I0(key1), .I1(rx_status2), .O(n874)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3521.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3522 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[35] ), 
            .O(n1247)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3522.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3523 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[34] ), 
            .O(n1251)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3523.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3524 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[33] ), 
            .O(n1254)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3524.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3525 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[39] ), 
            .O(n1261)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3525.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3526 (.I0(key2), .I1(\key2_counter[0] ), .O(n380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3526.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3527 (.I0(\key2_counter[0] ), .I1(\key2_counter[1] ), 
            .I2(\key2_counter[2] ), .I3(\key2_counter[3] ), .O(n2335)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3527.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3528 (.I0(n2335), .I1(\key2_counter[4] ), .I2(\key2_counter[5] ), 
            .I3(\key2_counter[6] ), .O(n2336)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf400 */ ;
    defparam LUT__3528.LUTMASK = 16'hf400;
    EFX_LUT4 LUT__3529 (.I0(\key2_counter[8] ), .I1(\key2_counter[9] ), 
            .O(n2337)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3529.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3530 (.I0(\key2_counter[10] ), .I1(\key2_counter[11] ), 
            .I2(\key2_counter[12] ), .I3(\key2_counter[13] ), .O(n2338)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3530.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3531 (.I0(\key2_counter[7] ), .I1(n2336), .I2(n2337), 
            .I3(n2338), .O(n2339)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1f00 */ ;
    defparam LUT__3531.LUTMASK = 16'h1f00;
    EFX_LUT4 LUT__3532 (.I0(key2), .I1(rx_status2), .I2(\key2_counter[14] ), 
            .I3(\key2_counter[15] ), .O(n2340)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3532.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3533 (.I0(\key1_counter[5] ), .I1(\key1_counter[7] ), 
            .I2(\key1_counter[6] ), .I3(\key1_counter[0]_2 ), .O(n2341)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3533.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3534 (.I0(\key1_counter[1] ), .I1(\key1_counter[2] ), 
            .I2(\key1_counter[4] ), .I3(\key1_counter[3] ), .O(n2342)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0100 */ ;
    defparam LUT__3534.LUTMASK = 16'h0100;
    EFX_LUT4 LUT__3535 (.I0(n2332), .I1(n2333), .I2(n2341), .I3(n2342), 
            .O(n2343)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3535.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3536 (.I0(n2340), .I1(n2339), .I2(n2343), .O(ceg_net83)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0d0d */ ;
    defparam LUT__3536.LUTMASK = 16'h0d0d;
    EFX_LUT4 LUT__3537 (.I0(\key2_counter[4] ), .I1(\key2_counter[3] ), 
            .I2(\key2_counter[0] ), .I3(\key2_counter[6] ), .O(n2344)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4000 */ ;
    defparam LUT__3537.LUTMASK = 16'h4000;
    EFX_LUT4 LUT__3538 (.I0(\key2_counter[1] ), .I1(\key2_counter[2] ), 
            .I2(\key2_counter[5] ), .I3(\key2_counter[7] ), .O(n2345)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3538.LUTMASK = 16'h0001;
    EFX_LUT4 LUT__3539 (.I0(\key2_counter[14] ), .I1(\key2_counter[15] ), 
            .I2(n2337), .O(n2346)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3539.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3540 (.I0(n2338), .I1(n2344), .I2(n2345), .I3(n2346), 
            .O(\equal_59/n31 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7fff */ ;
    defparam LUT__3540.LUTMASK = 16'h7fff;
    EFX_LUT4 LUT__3541 (.I0(n2343), .I1(rx_status2), .O(n875)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3541.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3542 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[38] ), 
            .O(n1272)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3542.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3543 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[36] ), 
            .O(n1277)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3543.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3544 (.I0(\r_mipi_rx_data_1P[31] ), .I1(\red_gain[1] ), 
            .O(n1280)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3544.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3545 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[37] ), 
            .O(n1282)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3545.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3546 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[36] ), 
            .O(n1288)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3546.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3547 (.I0(\key1_counter[0]_2 ), .I1(\key1_counter[1] ), 
            .O(n885)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3547.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3548 (.I0(\key1_counter[0]_2 ), .I1(\key1_counter[1] ), 
            .I2(\key1_counter[2] ), .O(n890)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3548.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3549 (.I0(\key1_counter[0]_2 ), .I1(\key1_counter[1] ), 
            .I2(\key1_counter[2] ), .I3(\key1_counter[3] ), .O(n895)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3549.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3550 (.I0(\key1_counter[0]_2 ), .I1(\key1_counter[1] ), 
            .I2(\key1_counter[2] ), .I3(\key1_counter[3] ), .O(n2347)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3550.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3551 (.I0(\key1_counter[4] ), .I1(n2347), .O(n900)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3551.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3552 (.I0(\key1_counter[4] ), .I1(n2347), .I2(\key1_counter[5] ), 
            .O(n905)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3552.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3553 (.I0(\key1_counter[4] ), .I1(\key1_counter[5] ), 
            .O(n2348)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3553.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3554 (.I0(n2347), .I1(n2348), .I2(\key1_counter[6] ), 
            .O(n910)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3554.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3555 (.I0(\key1_counter[6] ), .I1(n2347), .I2(n2348), 
            .I3(\key1_counter[7] ), .O(n915)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3555.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3556 (.I0(\key1_counter[6] ), .I1(\key1_counter[7] ), 
            .I2(n2347), .I3(n2348), .O(n2349)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3556.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3557 (.I0(\key1_counter[8] ), .I1(n2349), .O(n920)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3557.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3558 (.I0(\key1_counter[8] ), .I1(n2349), .I2(\key1_counter[9] ), 
            .O(n925)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3558.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3559 (.I0(\key1_counter[8] ), .I1(\key1_counter[9] ), 
            .I2(n2349), .I3(\key1_counter[10] ), .O(n930)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3559.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3560 (.I0(\key1_counter[8] ), .I1(\key1_counter[9] ), 
            .I2(\key1_counter[10] ), .O(n2350)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3560.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3561 (.I0(n2349), .I1(n2350), .O(n2351)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3561.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3562 (.I0(\key1_counter[11] ), .I1(n2351), .O(n935)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3562.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3563 (.I0(\key1_counter[11] ), .I1(n2351), .I2(\key1_counter[12] ), 
            .O(n940)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3563.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3564 (.I0(\key1_counter[11] ), .I1(\key1_counter[12] ), 
            .I2(n2349), .I3(n2350), .O(n2352)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3564.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3565 (.I0(\key1_counter[13] ), .I1(n2352), .O(n945)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3565.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3566 (.I0(\key1_counter[13] ), .I1(n2352), .I2(\key1_counter[14] ), 
            .O(n950)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3566.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3567 (.I0(\key1_counter[13] ), .I1(\key1_counter[14] ), 
            .I2(n2352), .I3(\key1_counter[15] ), .O(n955)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3567.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3568 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[35] ), 
            .O(n1309)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3568.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3569 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[34] ), 
            .O(n1312)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3569.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3570 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[33] ), 
            .O(n1315)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3570.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3571 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[32] ), 
            .O(n1318)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3571.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3572 (.I0(key2), .I1(\key2_counter[0] ), .I2(\key2_counter[1] ), 
            .O(n379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3572.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3573 (.I0(\key2_counter[0] ), .I1(\key2_counter[1] ), 
            .O(n2353)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3573.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3574 (.I0(key2), .I1(\key2_counter[2] ), .I2(n2353), 
            .O(n378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3574.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3575 (.I0(\key2_counter[2] ), .I1(n2353), .I2(key2), 
            .I3(\key2_counter[3] ), .O(n377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3575.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3576 (.I0(\key2_counter[0] ), .I1(\key2_counter[1] ), 
            .I2(\key2_counter[2] ), .I3(\key2_counter[3] ), .O(n2354)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3576.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3577 (.I0(key2), .I1(\key2_counter[4] ), .I2(n2354), 
            .O(n376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3577.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3578 (.I0(\key2_counter[4] ), .I1(n2354), .I2(key2), 
            .I3(\key2_counter[5] ), .O(n375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3578.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3579 (.I0(\key2_counter[4] ), .I1(\key2_counter[5] ), 
            .I2(n2354), .O(n2355)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3579.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3580 (.I0(key2), .I1(\key2_counter[6] ), .I2(n2355), 
            .O(n374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3580.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3581 (.I0(\key2_counter[6] ), .I1(n2355), .I2(key2), 
            .I3(\key2_counter[7] ), .O(n373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3581.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3582 (.I0(\key2_counter[6] ), .I1(\key2_counter[7] ), 
            .I2(n2355), .O(n2356)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3582.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3583 (.I0(key2), .I1(\key2_counter[8] ), .I2(n2356), 
            .O(n372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3583.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3584 (.I0(\key2_counter[8] ), .I1(n2356), .I2(key2), 
            .I3(\key2_counter[9] ), .O(n371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3584.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3585 (.I0(n2337), .I1(n2356), .I2(key2), .I3(\key2_counter[10] ), 
            .O(n370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3585.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3586 (.I0(\key2_counter[8] ), .I1(\key2_counter[9] ), 
            .I2(\key2_counter[10] ), .O(n2357)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3586.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3587 (.I0(n2356), .I1(n2357), .I2(key2), .I3(\key2_counter[11] ), 
            .O(n369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3587.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3588 (.I0(\key2_counter[6] ), .I1(\key2_counter[7] ), 
            .I2(\key2_counter[11] ), .I3(n2357), .O(n2358)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3588.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3589 (.I0(n2355), .I1(n2358), .I2(key2), .I3(\key2_counter[12] ), 
            .O(n368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3589.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3590 (.I0(\key2_counter[12] ), .I1(n2355), .I2(n2358), 
            .O(n2359)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3590.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3591 (.I0(key2), .I1(\key2_counter[13] ), .I2(n2359), 
            .O(n367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3591.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3592 (.I0(\key2_counter[12] ), .I1(\key2_counter[13] ), 
            .I2(n2355), .I3(n2358), .O(n2360)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3592.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3593 (.I0(key2), .I1(\key2_counter[14] ), .I2(n2360), 
            .O(n366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3593.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3594 (.I0(\key2_counter[14] ), .I1(n2360), .I2(key2), 
            .I3(\key2_counter[15] ), .O(n365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3594.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3595 (.I0(\red_gain[0] ), .I1(\red_gain[1] ), .O(n390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3595.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3596 (.I0(\red_gain[0] ), .I1(\red_gain[1] ), .I2(\red_gain[2] ), 
            .O(n389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3596.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3597 (.I0(\r_mipi_rx_data_1P[32] ), .I1(\red_gain[0] ), 
            .O(n1482)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3597.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3598 (.I0(\r_mipi_rx_data_1P[11] ), .I1(\red_gain[1] ), 
            .O(n1484)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3598.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3599 (.I0(\r_mipi_rx_data_1P[12] ), .I1(\red_gain[0] ), 
            .O(n1490)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3599.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3600 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[19] ), 
            .O(n1498)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3600.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3601 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[18] ), 
            .O(n1501)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3601.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3602 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[17] ), 
            .O(n1506)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3602.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3603 (.I0(n206), .I1(n413), .I2(\r_mipi_rx_data_1P[0] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/even_line_pix_0[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3603.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3604 (.I0(\inst_line_buf/r_mipi_rx_hsync_1P ), .I1(\inst_line_buf/r_mipi_rx_hsync_2P ), 
            .O(\inst_line_buf/n1283 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3604.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3605 (.I0(\inst_line_buf/r_mipi_rx_x_2P[0]_2 ), .I1(\inst_line_buf/n1283 ), 
            .O(\inst_line_buf/n1296 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3605.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3606 (.I0(\inst_line_buf/r_mipi_rx_valid_1P_2 ), .I1(\inst_line_buf/n1283 ), 
            .O(ceg_net98)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3606.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3607 (.I0(\inst_line_buf/r_mipi_tx_x_1P[0]_2 ), .I1(\inst_line_buf/r_mipi_tx_x_1P[1]_2 ), 
            .I2(\inst_line_buf/r_mipi_tx_x_1P[2]_2 ), .I3(\inst_line_buf/r_mipi_tx_x_1P[3]_2 ), 
            .O(n2361)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3607.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3608 (.I0(\inst_line_buf/r_mipi_tx_x_1P[5]_2 ), .I1(\inst_line_buf/r_mipi_tx_x_1P[9]_2 ), 
            .I2(\inst_line_buf/r_mipi_tx_x_1P[8]_2 ), .I3(\inst_line_buf/r_mipi_tx_x_1P[4]_2 ), 
            .O(n2362)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1000 */ ;
    defparam LUT__3608.LUTMASK = 16'h1000;
    EFX_LUT4 LUT__3609 (.I0(\inst_line_buf/r_mipi_tx_x_1P[6]_2 ), .I1(\inst_line_buf/r_mipi_tx_x_1P[7]_2 ), 
            .I2(n2361), .I3(n2362), .O(n2363)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3609.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3610 (.I0(\inst_line_buf/r_mipi_tx_x_inc_1P ), .I1(n2363), 
            .I2(\inst_line_buf/r_mipi_tx_en_1P ), .I3(\inst_line_buf/r_mipi_rx_full_1P_2 ), 
            .O(n2364)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h001f */ ;
    defparam LUT__3610.LUTMASK = 16'h001f;
    EFX_LUT4 LUT__3611 (.I0(n2363), .I1(\inst_line_buf/r_mipi_tx_x_inc_1P ), 
            .I2(\inst_line_buf/r_mipi_tx_en_1P ), .O(n2365)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4040 */ ;
    defparam LUT__3611.LUTMASK = 16'h4040;
    EFX_LUT4 LUT__3612 (.I0(n2365), .I1(n2364), .I2(\inst_line_buf/r_mipi_tx_x_1P[0]_2 ), 
            .O(\inst_line_buf/n1381 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3612.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3613 (.I0(\inst_line_buf/r_mipi_rx_full_1P_2 ), .I1(\inst_line_buf/n1283 ), 
            .O(ceg_net101)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3613.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3614 (.I0(\inst_line_buf/r_mipi_tx_en_1P ), .I1(n2363), 
            .O(\inst_line_buf/n2531 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3614.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3615 (.I0(\inst_line_buf/r_mipi_rx_full_1P_2 ), .I1(\inst_line_buf/n2531 ), 
            .O(ceg_net104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3615.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3616 (.I0(\inst_line_buf/r_mipi_tx_b_1P[0] ), .I1(\inst_line_buf/r_mipi_tx_b_1P[2] ), 
            .I2(\inst_line_buf/r_mipi_tx_b_1P[1] ), .I3(\inst_line_buf/r_mipi_tx_en_1P ), 
            .O(\inst_line_buf/n1387 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hef00 */ ;
    defparam LUT__3616.LUTMASK = 16'hef00;
    EFX_LUT4 LUT__3617 (.I0(n2363), .I1(\inst_line_buf/n1387 ), .O(n2366)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3617.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3618 (.I0(\inst_line_buf/r_mipi_tx_b_1P[0] ), .I1(n2366), 
            .O(\inst_line_buf/n1385 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3618.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3619 (.I0(\inst_line_buf/r_mipi_rx_full_1P_2 ), .I1(\inst_line_buf/r_mipi_tx_en_1P ), 
            .O(ceg_net140)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1111 */ ;
    defparam LUT__3619.LUTMASK = 16'h1111;
    EFX_LUT4 LUT__3620 (.I0(\inst_line_buf/r_mipi_tx_data_5P[60] ), .I1(\inst_line_buf/r_mipi_tx_data_4P[0] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1510 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hacac */ ;
    defparam LUT__3620.LUTMASK = 16'hacac;
    EFX_LUT4 LUT__3621 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[16] ), 
            .O(n1533)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3621.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3622 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[31] ), 
            .O(n1548)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3622.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3623 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[32] ), 
            .O(n1550)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3623.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3624 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[11] ), 
            .O(n1553)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3624.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3625 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[12] ), 
            .O(n1555)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3625.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3626 (.I0(n206), .I1(n223), .I2(\r_mipi_rx_data_1P[1] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3626.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3627 (.I0(n206), .I1(n221), .I2(\r_mipi_rx_data_1P[2] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3627.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3628 (.I0(n206), .I1(n219), .I2(\r_mipi_rx_data_1P[3] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3628.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3629 (.I0(n206), .I1(n217), .I2(\r_mipi_rx_data_1P[4] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3629.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3630 (.I0(n206), .I1(n215), .I2(\r_mipi_rx_data_1P[5] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3630.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3631 (.I0(n206), .I1(n213), .I2(\r_mipi_rx_data_1P[6] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3631.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3632 (.I0(n206), .I1(n211), .I2(\r_mipi_rx_data_1P[7] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3632.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3633 (.I0(n206), .I1(n209), .I2(\r_mipi_rx_data_1P[8] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3633.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3634 (.I0(n206), .I1(n207), .I2(\r_mipi_rx_data_1P[9] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_0[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3634.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3635 (.I0(n423), .I1(n355), .I2(\red_gain[2] ), .O(n2367)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3635.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3636 (.I0(n354), .I1(n883), .I2(\red_gain[2] ), .O(n2368)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3636.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3637 (.I0(n247), .I1(n407), .I2(\r_mipi_rx_data_1P[10] ), 
            .I3(\green_gain[2] ), .O(n2369)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3637.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3638 (.I0(n2368), .I1(n2367), .I2(n2369), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[10] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3638.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3639 (.I0(n943), .I1(n900_2), .I2(\red_gain[2] ), .O(n2370)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3639.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3640 (.I0(n247), .I1(n264), .I2(\r_mipi_rx_data_1P[11] ), 
            .I3(\green_gain[2] ), .O(n2371)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3640.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3641 (.I0(n2368), .I1(n2370), .I2(n2371), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[11] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3641.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3642 (.I0(n941), .I1(n898), .I2(\red_gain[2] ), .O(n2372)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3642.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3643 (.I0(n247), .I1(n262), .I2(\r_mipi_rx_data_1P[12] ), 
            .I3(\green_gain[2] ), .O(n2373)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3643.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3644 (.I0(n2368), .I1(n2372), .I2(n2373), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[12] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3644.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3645 (.I0(n939), .I1(n896), .I2(\red_gain[2] ), .O(n2374)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3645.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3646 (.I0(n247), .I1(n260), .I2(\r_mipi_rx_data_1P[13] ), 
            .I3(\green_gain[2] ), .O(n2375)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3646.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3647 (.I0(n2368), .I1(n2374), .I2(n2375), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[13] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3647.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3648 (.I0(n394), .I1(n894), .I2(\red_gain[2] ), .O(n2376)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3648.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3649 (.I0(n247), .I1(n258), .I2(\r_mipi_rx_data_1P[14] ), 
            .I3(\green_gain[2] ), .O(n2377)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3649.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3650 (.I0(n2368), .I1(n2376), .I2(n2377), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[14] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3650.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3651 (.I0(n371_2), .I1(n892), .I2(\red_gain[2] ), .O(n2378)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3651.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3652 (.I0(n247), .I1(n256), .I2(\r_mipi_rx_data_1P[15] ), 
            .I3(\green_gain[2] ), .O(n2379)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3652.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3653 (.I0(n2368), .I1(n2378), .I2(n2379), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[15] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3653.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3654 (.I0(n367_2), .I1(n890_2), .I2(\red_gain[2] ), 
            .O(n2380)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3654.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3655 (.I0(n247), .I1(n254), .I2(\r_mipi_rx_data_1P[16] ), 
            .I3(\green_gain[2] ), .O(n2381)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3655.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3656 (.I0(n2368), .I1(n2380), .I2(n2381), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[16] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3656.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3657 (.I0(n365_2), .I1(n888), .I2(\red_gain[2] ), .O(n2382)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3657.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3658 (.I0(n247), .I1(n252), .I2(\r_mipi_rx_data_1P[17] ), 
            .I3(\green_gain[2] ), .O(n2383)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3658.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3659 (.I0(n2368), .I1(n2382), .I2(n2383), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[17] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3659.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3660 (.I0(n361), .I1(n886), .I2(\red_gain[2] ), .O(n2384)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3660.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3661 (.I0(n247), .I1(n250), .I2(\r_mipi_rx_data_1P[18] ), 
            .I3(\green_gain[2] ), .O(n2385)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3661.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3662 (.I0(n2368), .I1(n2384), .I2(n2385), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[18] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3662.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3663 (.I0(n359), .I1(n884), .I2(\red_gain[2] ), .O(n2386)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3663.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3664 (.I0(n247), .I1(n248), .I2(\r_mipi_rx_data_1P[19] ), 
            .I3(\green_gain[2] ), .O(n2387)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3664.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3665 (.I0(n2368), .I1(n2386), .I2(n2387), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[19] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3665.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3666 (.I0(n401), .I1(n1034), .I2(\r_mipi_rx_data_1P[20] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/even_line_pix_2[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3666.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3667 (.I0(n1034), .I1(n1051), .I2(\r_mipi_rx_data_1P[21] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[1] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3667.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3668 (.I0(n1034), .I1(n1049), .I2(\r_mipi_rx_data_1P[22] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[2] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3668.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3669 (.I0(n1034), .I1(n1047), .I2(\r_mipi_rx_data_1P[23] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[3] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3669.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3670 (.I0(n1034), .I1(n1045), .I2(\r_mipi_rx_data_1P[24] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[4] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3670.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3671 (.I0(n1034), .I1(n1043), .I2(\r_mipi_rx_data_1P[25] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[5] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3671.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3672 (.I0(n1034), .I1(n1041), .I2(\r_mipi_rx_data_1P[26] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[6] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3672.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3673 (.I0(n1034), .I1(n1039), .I2(\r_mipi_rx_data_1P[27] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[7] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3673.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3674 (.I0(n1034), .I1(n1037), .I2(\r_mipi_rx_data_1P[28] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[8] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3674.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3675 (.I0(n1034), .I1(n1035), .I2(\r_mipi_rx_data_1P[29] ), 
            .I3(\green_gain[2] ), .O(\inst_line_buf/odd_line_pix_2[9] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3675.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3676 (.I0(n417), .I1(n348), .I2(\red_gain[2] ), .O(n2388)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3676.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3677 (.I0(n1081), .I1(n920_2), .I2(\red_gain[2] ), .O(n2389)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3677.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3678 (.I0(n363), .I1(n845), .I2(\r_mipi_rx_data_1P[30] ), 
            .I3(\green_gain[2] ), .O(n2390)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3678.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3679 (.I0(n2389), .I1(n2388), .I2(n2390), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[30] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3679.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3680 (.I0(n937), .I1(n155), .I2(\red_gain[2] ), .O(n2391)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3680.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3681 (.I0(n845), .I1(n862), .I2(\r_mipi_rx_data_1P[31] ), 
            .I3(\green_gain[2] ), .O(n2392)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3681.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3682 (.I0(n2389), .I1(n2391), .I2(n2392), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[31] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3682.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3683 (.I0(n935_2), .I1(n153), .I2(\red_gain[2] ), .O(n2393)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3683.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3684 (.I0(n845), .I1(n860), .I2(\r_mipi_rx_data_1P[32] ), 
            .I3(\green_gain[2] ), .O(n2394)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3684.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3685 (.I0(n2389), .I1(n2393), .I2(n2394), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[32] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3685.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3686 (.I0(n933), .I1(n150), .I2(\red_gain[2] ), .O(n2395)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3686.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3687 (.I0(n845), .I1(n858), .I2(\r_mipi_rx_data_1P[33] ), 
            .I3(\green_gain[2] ), .O(n2396)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3687.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3688 (.I0(n2389), .I1(n2395), .I2(n2396), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[33] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3688.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3689 (.I0(n931), .I1(n171_2), .I2(\red_gain[2] ), .O(n2397)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h5353 */ ;
    defparam LUT__3689.LUTMASK = 16'h5353;
    EFX_LUT4 LUT__3690 (.I0(n845), .I1(n856), .I2(\r_mipi_rx_data_1P[34] ), 
            .I3(\green_gain[2] ), .O(n2398)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3690.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3691 (.I0(n2389), .I1(n2397), .I2(n2398), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[34] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3691.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3692 (.I0(n1090_2), .I1(n929), .I2(\red_gain[2] ), .O(n2399)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3692.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3693 (.I0(n845), .I1(n854), .I2(\r_mipi_rx_data_1P[35] ), 
            .I3(\green_gain[2] ), .O(n2400)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3693.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3694 (.I0(n2389), .I1(n2399), .I2(n2400), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[35] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3694.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3695 (.I0(n1088), .I1(n927), .I2(\red_gain[2] ), .O(n2401)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3695.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3696 (.I0(n845), .I1(n852), .I2(\r_mipi_rx_data_1P[36] ), 
            .I3(\green_gain[2] ), .O(n2402)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3696.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3697 (.I0(n2389), .I1(n2401), .I2(n2402), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[36] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3697.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3698 (.I0(n1086), .I1(n925_2), .I2(\red_gain[2] ), .O(n2403)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3698.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3699 (.I0(n845), .I1(n850), .I2(\r_mipi_rx_data_1P[37] ), 
            .I3(\green_gain[2] ), .O(n2404)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3699.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3700 (.I0(n2389), .I1(n2403), .I2(n2404), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[37] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3700.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3701 (.I0(n1084), .I1(n923), .I2(\red_gain[2] ), .O(n2405)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3701.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3702 (.I0(n845), .I1(n848), .I2(\r_mipi_rx_data_1P[38] ), 
            .I3(\green_gain[2] ), .O(n2406)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3702.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3703 (.I0(n2389), .I1(n2405), .I2(n2406), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[38] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3703.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3704 (.I0(n1082), .I1(n921), .I2(\red_gain[2] ), .O(n2407)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h3535 */ ;
    defparam LUT__3704.LUTMASK = 16'h3535;
    EFX_LUT4 LUT__3705 (.I0(n845), .I1(n846), .I2(\r_mipi_rx_data_1P[39] ), 
            .I3(\green_gain[2] ), .O(n2408)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hf0ee */ ;
    defparam LUT__3705.LUTMASK = 16'hf0ee;
    EFX_LUT4 LUT__3706 (.I0(n2389), .I1(n2407), .I2(n2408), .I3(\inst_line_buf/r_mipi_rx_x_2P[10]_2 ), 
            .O(\inst_line_buf/mipi_inst1_DATA_filtered[39] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h77f0 */ ;
    defparam LUT__3706.LUTMASK = 16'h77f0;
    EFX_LUT4 LUT__3707 (.I0(\inst_line_buf/n1283 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[0]_2 ), 
            .I2(\inst_line_buf/r_mipi_rx_x_2P[1]_2 ), .O(\inst_line_buf/n1295 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3707.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3708 (.I0(\inst_line_buf/r_mipi_rx_x_2P[0]_2 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[1]_2 ), 
            .O(n2409)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3708.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3709 (.I0(\inst_line_buf/n1283 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[2]_2 ), 
            .I2(n2409), .O(\inst_line_buf/n1294 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3709.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3710 (.I0(\inst_line_buf/r_mipi_rx_x_2P[2]_2 ), .I1(n2409), 
            .I2(\inst_line_buf/n1283 ), .I3(\inst_line_buf/r_mipi_rx_x_2P[3]_2 ), 
            .O(\inst_line_buf/n1293 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3710.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3711 (.I0(\inst_line_buf/r_mipi_rx_x_2P[0]_2 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[1]_2 ), 
            .I2(\inst_line_buf/r_mipi_rx_x_2P[2]_2 ), .I3(\inst_line_buf/r_mipi_rx_x_2P[3]_2 ), 
            .O(n2410)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3711.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3712 (.I0(\inst_line_buf/n1283 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[4]_2 ), 
            .I2(n2410), .O(\inst_line_buf/n1292 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3712.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3713 (.I0(\inst_line_buf/r_mipi_rx_x_2P[4]_2 ), .I1(n2410), 
            .I2(\inst_line_buf/n1283 ), .I3(\inst_line_buf/r_mipi_rx_x_2P[5]_2 ), 
            .O(\inst_line_buf/n1291 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3713.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3714 (.I0(\inst_line_buf/r_mipi_rx_x_2P[4]_2 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[5]_2 ), 
            .I2(n2410), .O(n2411)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3714.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3715 (.I0(\inst_line_buf/n1283 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[6]_2 ), 
            .I2(n2411), .O(\inst_line_buf/n1290 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3715.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3716 (.I0(\inst_line_buf/r_mipi_rx_x_2P[6]_2 ), .I1(n2411), 
            .I2(\inst_line_buf/n1283 ), .I3(\inst_line_buf/r_mipi_rx_x_2P[7]_2 ), 
            .O(\inst_line_buf/n1289 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3716.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3717 (.I0(\inst_line_buf/r_mipi_rx_x_2P[6]_2 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[7]_2 ), 
            .I2(n2411), .O(n2412)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8080 */ ;
    defparam LUT__3717.LUTMASK = 16'h8080;
    EFX_LUT4 LUT__3718 (.I0(\inst_line_buf/n1283 ), .I1(\inst_line_buf/r_mipi_rx_x_2P[8]_2 ), 
            .I2(n2412), .O(\inst_line_buf/n1288 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h1414 */ ;
    defparam LUT__3718.LUTMASK = 16'h1414;
    EFX_LUT4 LUT__3719 (.I0(\inst_line_buf/r_mipi_rx_x_2P[8]_2 ), .I1(n2412), 
            .I2(\inst_line_buf/n1283 ), .I3(\inst_line_buf/r_mipi_rx_x_2P[9]_2 ), 
            .O(\inst_line_buf/n1287 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0708 */ ;
    defparam LUT__3719.LUTMASK = 16'h0708;
    EFX_LUT4 LUT__3720 (.I0(n2364), .I1(\inst_line_buf/r_mipi_tx_x_1P[0]_2 ), 
            .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[1]_2 ), .O(\inst_line_buf/n1380 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3720.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3721 (.I0(\inst_line_buf/r_mipi_tx_x_1P[0]_2 ), .I1(\inst_line_buf/r_mipi_tx_x_1P[1]_2 ), 
            .O(n2413)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3721.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3722 (.I0(n2364), .I1(n2413), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[2]_2 ), 
            .O(\inst_line_buf/n1379 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3722.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3723 (.I0(\inst_line_buf/r_mipi_tx_x_1P[2]_2 ), .I1(n2413), 
            .O(n2414)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3723.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3724 (.I0(n2364), .I1(n2414), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[3]_2 ), 
            .O(\inst_line_buf/n1378 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3724.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3725 (.I0(n2364), .I1(n2361), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[4]_2 ), 
            .O(\inst_line_buf/n1377 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3725.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3726 (.I0(\inst_line_buf/r_mipi_tx_x_1P[4]_2 ), .I1(n2361), 
            .O(n2415)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3726.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3727 (.I0(n2364), .I1(n2415), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[5]_2 ), 
            .O(\inst_line_buf/n1376 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3727.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3728 (.I0(\inst_line_buf/r_mipi_tx_x_1P[4]_2 ), .I1(\inst_line_buf/r_mipi_tx_x_1P[5]_2 ), 
            .O(n2416)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3728.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3729 (.I0(n2361), .I1(n2416), .O(n2417)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3729.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3730 (.I0(n2364), .I1(n2417), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[6]_2 ), 
            .O(\inst_line_buf/n1375 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3730.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3731 (.I0(\inst_line_buf/r_mipi_tx_x_1P[6]_2 ), .I1(n2417), 
            .O(n2418)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3731.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3732 (.I0(n2364), .I1(n2418), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[7]_2 ), 
            .O(\inst_line_buf/n1374 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3732.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3733 (.I0(\inst_line_buf/r_mipi_tx_x_1P[6]_2 ), .I1(\inst_line_buf/r_mipi_tx_x_1P[7]_2 ), 
            .I2(n2361), .I3(n2416), .O(n2419)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3733.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3734 (.I0(n2364), .I1(n2419), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[8]_2 ), 
            .O(\inst_line_buf/n1373 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3734.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3735 (.I0(\inst_line_buf/r_mipi_tx_x_1P[6]_2 ), .I1(\inst_line_buf/r_mipi_tx_x_1P[7]_2 ), 
            .I2(\inst_line_buf/r_mipi_tx_x_1P[8]_2 ), .I3(n2417), .O(n2420)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3735.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3736 (.I0(n2364), .I1(n2420), .I2(n2365), .I3(\inst_line_buf/r_mipi_tx_x_1P[9]_2 ), 
            .O(\inst_line_buf/n1372 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbac0 */ ;
    defparam LUT__3736.LUTMASK = 16'hbac0;
    EFX_LUT4 LUT__3737 (.I0(\inst_line_buf/r_mipi_tx_b_1P[0] ), .I1(\inst_line_buf/r_mipi_tx_b_1P[1] ), 
            .I2(n2366), .O(\inst_line_buf/n1384 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6060 */ ;
    defparam LUT__3737.LUTMASK = 16'h6060;
    EFX_LUT4 LUT__3738 (.I0(\inst_line_buf/r_mipi_tx_b_1P[0] ), .I1(\inst_line_buf/r_mipi_tx_b_1P[1] ), 
            .I2(\inst_line_buf/r_mipi_tx_b_1P[2] ), .I3(n2366), .O(\inst_line_buf/n1383 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7800 */ ;
    defparam LUT__3738.LUTMASK = 16'h7800;
    EFX_LUT4 LUT__3739 (.I0(\inst_line_buf/r_mipi_tx_data_4P[1] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[61] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1509 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3739.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3740 (.I0(\inst_line_buf/r_mipi_tx_data_4P[2] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[62] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1508 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3740.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3741 (.I0(\inst_line_buf/r_mipi_tx_data_4P[3] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[63] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1507 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3741.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3742 (.I0(\inst_line_buf/r_mipi_tx_data_4P[4] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[64] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1506 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3742.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3743 (.I0(\inst_line_buf/r_mipi_tx_data_4P[5] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[65] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1505 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3743.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3744 (.I0(\inst_line_buf/r_mipi_tx_data_4P[6] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[66] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1504 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3744.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3745 (.I0(\inst_line_buf/r_mipi_tx_data_4P[7] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[67] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1503 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3745.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3746 (.I0(\inst_line_buf/r_mipi_tx_data_4P[8] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[68] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1502 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3746.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3747 (.I0(\inst_line_buf/r_mipi_tx_data_4P[9] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[69] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1501 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3747.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3748 (.I0(\inst_line_buf/r_mipi_tx_data_4P[10] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[70] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1500 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3748.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3749 (.I0(\inst_line_buf/r_mipi_tx_data_4P[11] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[71] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1499 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3749.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3750 (.I0(\inst_line_buf/r_mipi_tx_data_4P[12] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[72] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1498 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3750.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3751 (.I0(\inst_line_buf/r_mipi_tx_data_4P[13] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[73] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1497 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3751.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3752 (.I0(\inst_line_buf/r_mipi_tx_data_4P[14] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[74] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1496 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3752.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3753 (.I0(\inst_line_buf/r_mipi_tx_data_4P[15] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[75] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1495 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3753.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3754 (.I0(\inst_line_buf/r_mipi_tx_data_4P[16] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[76] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1494 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3754.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3755 (.I0(\inst_line_buf/r_mipi_tx_data_4P[17] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[77] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1493 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3755.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3756 (.I0(\inst_line_buf/r_mipi_tx_data_4P[18] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[78] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1492 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3756.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3757 (.I0(\inst_line_buf/r_mipi_tx_data_4P[19] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[79] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1491 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3757.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3758 (.I0(\inst_line_buf/r_mipi_tx_data_4P[20] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[80] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1490 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3758.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3759 (.I0(\inst_line_buf/r_mipi_tx_data_4P[21] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[81] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1489 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3759.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3760 (.I0(\inst_line_buf/r_mipi_tx_data_4P[22] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[82] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1488 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3760.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3761 (.I0(\inst_line_buf/r_mipi_tx_data_4P[23] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[83] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1487 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3761.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3762 (.I0(\inst_line_buf/r_mipi_tx_data_4P[24] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[84] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1486 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3762.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3763 (.I0(\inst_line_buf/r_mipi_tx_data_4P[25] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[85] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1485 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3763.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3764 (.I0(\inst_line_buf/r_mipi_tx_data_4P[26] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[86] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1484 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3764.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3765 (.I0(\inst_line_buf/r_mipi_tx_data_4P[27] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[87] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1483 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3765.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3766 (.I0(\inst_line_buf/r_mipi_tx_data_4P[28] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[88] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1482 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3766.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3767 (.I0(\inst_line_buf/r_mipi_tx_data_4P[29] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[89] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1481 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3767.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3768 (.I0(\inst_line_buf/r_mipi_tx_data_4P[30] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[90] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1480 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3768.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3769 (.I0(\inst_line_buf/r_mipi_tx_data_4P[31] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[91] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1479 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3769.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3770 (.I0(\inst_line_buf/r_mipi_tx_data_4P[32] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[92] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1478 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3770.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3771 (.I0(\inst_line_buf/r_mipi_tx_data_4P[33] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[93] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1477 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3771.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3772 (.I0(\inst_line_buf/r_mipi_tx_data_4P[34] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[94] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1476 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3772.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3773 (.I0(\inst_line_buf/r_mipi_tx_data_4P[35] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[95] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1475 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3773.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3774 (.I0(\inst_line_buf/r_mipi_tx_data_4P[36] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[96] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1474 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3774.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3775 (.I0(\inst_line_buf/r_mipi_tx_data_4P[37] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[97] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1473 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3775.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3776 (.I0(\inst_line_buf/r_mipi_tx_data_4P[38] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[98] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1472 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3776.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3777 (.I0(\inst_line_buf/r_mipi_tx_data_4P[39] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[99] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1471 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3777.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3778 (.I0(\inst_line_buf/r_mipi_tx_data_4P[40] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[100] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1470 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3778.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3779 (.I0(\inst_line_buf/r_mipi_tx_data_4P[41] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[101] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1469 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3779.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3780 (.I0(\inst_line_buf/r_mipi_tx_data_4P[42] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[102] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1468 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3780.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3781 (.I0(\inst_line_buf/r_mipi_tx_data_4P[43] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[103] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1467 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3781.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3782 (.I0(\inst_line_buf/r_mipi_tx_data_4P[44] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[104] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1466 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3782.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3783 (.I0(\inst_line_buf/r_mipi_tx_data_4P[45] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[105] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1465 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3783.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3784 (.I0(\inst_line_buf/r_mipi_tx_data_4P[46] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[106] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1464 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3784.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3785 (.I0(\inst_line_buf/r_mipi_tx_data_4P[47] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[107] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1463 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3785.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3786 (.I0(\inst_line_buf/r_mipi_tx_data_4P[48] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[108] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1462 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3786.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3787 (.I0(\inst_line_buf/r_mipi_tx_data_4P[49] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[109] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1461 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3787.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3788 (.I0(\inst_line_buf/r_mipi_tx_data_4P[50] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[110] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1460 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3788.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3789 (.I0(\inst_line_buf/r_mipi_tx_data_4P[51] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[111] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1459 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3789.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3790 (.I0(\inst_line_buf/r_mipi_tx_data_4P[52] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[112] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1458 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3790.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3791 (.I0(\inst_line_buf/r_mipi_tx_data_4P[53] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[113] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1457 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3791.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3792 (.I0(\inst_line_buf/r_mipi_tx_data_4P[54] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[114] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1456 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3792.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3793 (.I0(\inst_line_buf/r_mipi_tx_data_4P[55] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[115] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1455 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3793.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3794 (.I0(\inst_line_buf/r_mipi_tx_data_4P[56] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[116] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1454 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3794.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3795 (.I0(\inst_line_buf/r_mipi_tx_data_4P[57] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[117] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1453 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3795.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3796 (.I0(\inst_line_buf/r_mipi_tx_data_4P[58] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[118] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1452 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3796.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3797 (.I0(\inst_line_buf/r_mipi_tx_data_4P[59] ), .I1(\inst_line_buf/r_mipi_tx_data_5P[119] ), 
            .I2(mipi_inst2_VALID), .O(\inst_line_buf/n1451 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3797.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3798 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[60] ), 
            .O(\inst_line_buf/n1450 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3798.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3799 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[61] ), 
            .O(\inst_line_buf/n1449 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3799.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3800 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[62] ), 
            .O(\inst_line_buf/n1448 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3800.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3801 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[63] ), 
            .O(\inst_line_buf/n1447 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3801.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3802 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[64] ), 
            .O(\inst_line_buf/n1446 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3802.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3803 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[65] ), 
            .O(\inst_line_buf/n1445 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3803.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3804 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[66] ), 
            .O(\inst_line_buf/n1444 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3804.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3805 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[67] ), 
            .O(\inst_line_buf/n1443 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3805.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3806 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[68] ), 
            .O(\inst_line_buf/n1442 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3806.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3807 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[69] ), 
            .O(\inst_line_buf/n1441 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3807.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3808 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[70] ), 
            .O(\inst_line_buf/n1440 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3808.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3809 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[71] ), 
            .O(\inst_line_buf/n1439 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3809.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3810 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[72] ), 
            .O(\inst_line_buf/n1438 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3810.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3811 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[73] ), 
            .O(\inst_line_buf/n1437 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3811.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3812 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[74] ), 
            .O(\inst_line_buf/n1436 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3812.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3813 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[75] ), 
            .O(\inst_line_buf/n1435 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3813.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3814 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[76] ), 
            .O(\inst_line_buf/n1434 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3814.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3815 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[77] ), 
            .O(\inst_line_buf/n1433 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3815.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3816 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[78] ), 
            .O(\inst_line_buf/n1432 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3816.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3817 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[79] ), 
            .O(\inst_line_buf/n1431 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3817.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3818 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[80] ), 
            .O(\inst_line_buf/n1430 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3818.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3819 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[81] ), 
            .O(\inst_line_buf/n1429 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3819.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3820 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[82] ), 
            .O(\inst_line_buf/n1428 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3820.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3821 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[83] ), 
            .O(\inst_line_buf/n1427 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3821.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3822 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[84] ), 
            .O(\inst_line_buf/n1426 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3822.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3823 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[85] ), 
            .O(\inst_line_buf/n1425 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3823.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3824 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[86] ), 
            .O(\inst_line_buf/n1424 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3824.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3825 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[87] ), 
            .O(\inst_line_buf/n1423 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3825.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3826 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[88] ), 
            .O(\inst_line_buf/n1422 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3826.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3827 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[89] ), 
            .O(\inst_line_buf/n1421 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3827.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3828 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[90] ), 
            .O(\inst_line_buf/n1420 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3828.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3829 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[91] ), 
            .O(\inst_line_buf/n1419 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3829.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3830 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[92] ), 
            .O(\inst_line_buf/n1418 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3830.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3831 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[93] ), 
            .O(\inst_line_buf/n1417 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3831.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3832 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[94] ), 
            .O(\inst_line_buf/n1416 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3832.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3833 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[95] ), 
            .O(\inst_line_buf/n1415 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3833.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3834 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[96] ), 
            .O(\inst_line_buf/n1414 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3834.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3835 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[97] ), 
            .O(\inst_line_buf/n1413 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3835.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3836 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[98] ), 
            .O(\inst_line_buf/n1412 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3836.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3837 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[99] ), 
            .O(\inst_line_buf/n1411 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3837.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3838 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[100] ), 
            .O(\inst_line_buf/n1410 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3838.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3839 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[101] ), 
            .O(\inst_line_buf/n1409 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3839.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3840 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[102] ), 
            .O(\inst_line_buf/n1408 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3840.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3841 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[103] ), 
            .O(\inst_line_buf/n1407 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3841.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3842 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[104] ), 
            .O(\inst_line_buf/n1406 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3842.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3843 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[105] ), 
            .O(\inst_line_buf/n1405 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3843.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3844 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[106] ), 
            .O(\inst_line_buf/n1404 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3844.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3845 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[107] ), 
            .O(\inst_line_buf/n1403 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3845.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3846 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[108] ), 
            .O(\inst_line_buf/n1402 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3846.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3847 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[109] ), 
            .O(\inst_line_buf/n1401 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3847.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3848 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[110] ), 
            .O(\inst_line_buf/n1400 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3848.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3849 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[111] ), 
            .O(\inst_line_buf/n1399 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3849.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3850 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[112] ), 
            .O(\inst_line_buf/n1398 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3850.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3851 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[113] ), 
            .O(\inst_line_buf/n1397 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3851.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3852 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[114] ), 
            .O(\inst_line_buf/n1396 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3852.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3853 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[115] ), 
            .O(\inst_line_buf/n1395 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3853.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3854 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[116] ), 
            .O(\inst_line_buf/n1394 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3854.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3855 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[117] ), 
            .O(\inst_line_buf/n1393 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3855.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3856 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[118] ), 
            .O(\inst_line_buf/n1392 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3856.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3857 (.I0(mipi_inst2_VALID), .I1(\inst_line_buf/r_mipi_tx_data_4P[119] ), 
            .O(\inst_line_buf/n1391 )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3857.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3858 (.I0(r_rden_1P_2), .I1(\r_raddr_1P[12]_2 ), .O(n1502)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3858.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3859 (.I0(\r_mipi_rx_data_1P[19] ), .I1(\red_gain[0] ), 
            .O(n2071)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3859.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3860 (.I0(\r_mipi_rx_data_1P[18] ), .I1(\red_gain[0] ), 
            .O(n2074)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3860.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3861 (.I0(\r_mipi_rx_data_1P[17] ), .I1(\red_gain[0] ), 
            .O(n2077)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3861.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3862 (.I0(\r_mipi_rx_data_1P[16] ), .I1(\red_gain[0] ), 
            .O(n2080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3862.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3863 (.I0(\r_mipi_rx_data_1P[15] ), .I1(\red_gain[0] ), 
            .O(n2083)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3863.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3864 (.I0(\r_mipi_rx_data_1P[14] ), .I1(\red_gain[0] ), 
            .O(n2086)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3864.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3865 (.I0(\r_mipi_rx_data_1P[13] ), .I1(\red_gain[0] ), 
            .O(n2089)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3865.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3866 (.I0(\r_mipi_rx_data_1P[19] ), .I1(\red_gain[1] ), 
            .O(n2092)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3866.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3867 (.I0(\r_mipi_rx_data_1P[18] ), .I1(\red_gain[1] ), 
            .O(n2094)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3867.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3868 (.I0(\r_mipi_rx_data_1P[17] ), .I1(\red_gain[1] ), 
            .O(n2096)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3868.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3869 (.I0(\r_mipi_rx_data_1P[16] ), .I1(\red_gain[1] ), 
            .O(n2098)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3869.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3870 (.I0(\r_mipi_rx_data_1P[15] ), .I1(\red_gain[1] ), 
            .O(n2100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3870.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3871 (.I0(\r_mipi_rx_data_1P[14] ), .I1(\red_gain[1] ), 
            .O(n2102)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3871.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3872 (.I0(\r_mipi_rx_data_1P[13] ), .I1(\red_gain[1] ), 
            .O(n2104)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3872.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3873 (.I0(\r_mipi_rx_data_1P[12] ), .I1(\red_gain[1] ), 
            .O(n2106)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3873.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3874 (.I0(\r_mipi_rx_data_1P[39] ), .I1(\red_gain[0] ), 
            .O(n2115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3874.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3875 (.I0(\r_mipi_rx_data_1P[38] ), .I1(\red_gain[0] ), 
            .O(n2118)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3875.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3876 (.I0(\r_mipi_rx_data_1P[37] ), .I1(\red_gain[0] ), 
            .O(n2121)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3876.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3877 (.I0(\r_mipi_rx_data_1P[36] ), .I1(\red_gain[0] ), 
            .O(n2124)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3877.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3878 (.I0(\r_mipi_rx_data_1P[35] ), .I1(\red_gain[0] ), 
            .O(n2127)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3878.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3879 (.I0(\r_mipi_rx_data_1P[34] ), .I1(\red_gain[0] ), 
            .O(n2130)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3879.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3880 (.I0(\r_mipi_rx_data_1P[33] ), .I1(\red_gain[0] ), 
            .O(n2133)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3880.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3881 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[15] ), 
            .O(n2136)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3881.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3882 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[14] ), 
            .O(n2139)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3882.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3883 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[13] ), 
            .O(n2142)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3883.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3884 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[19] ), 
            .O(n2146)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3884.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3885 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[18] ), 
            .O(n2148)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3885.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3886 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[17] ), 
            .O(n2150)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3886.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3887 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[16] ), 
            .O(n2152)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3887.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3888 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[15] ), 
            .O(n2154)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3888.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3889 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[14] ), 
            .O(n2156)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3889.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3890 (.I0(\r_mipi_rx_data_1P[39] ), .I1(\red_gain[1] ), 
            .O(n2159)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3890.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3891 (.I0(\r_mipi_rx_data_1P[38] ), .I1(\red_gain[1] ), 
            .O(n2161)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3891.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3892 (.I0(\r_mipi_rx_data_1P[37] ), .I1(\red_gain[1] ), 
            .O(n2163)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3892.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3893 (.I0(\r_mipi_rx_data_1P[36] ), .I1(\red_gain[1] ), 
            .O(n2165)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3893.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3894 (.I0(\r_mipi_rx_data_1P[35] ), .I1(\red_gain[1] ), 
            .O(n2167)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3894.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3895 (.I0(\r_mipi_rx_data_1P[34] ), .I1(\red_gain[1] ), 
            .O(n2169)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3895.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3896 (.I0(\r_mipi_rx_data_1P[33] ), .I1(\red_gain[1] ), 
            .O(n2171)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3896.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3897 (.I0(\r_mipi_rx_data_1P[32] ), .I1(\red_gain[1] ), 
            .O(n2173)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3897.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3898 (.I0(\r_raddr_1P[0]_2 ), .I1(\r_raddr_1P[1]_2 ), 
            .O(n1060)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3898.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3899 (.I0(\r_raddr_1P[0]_2 ), .I1(\r_raddr_1P[1]_2 ), 
            .I2(\r_raddr_1P[2]_2 ), .O(n1065)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3899.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3900 (.I0(\r_raddr_1P[0]_2 ), .I1(\r_raddr_1P[1]_2 ), 
            .I2(\r_raddr_1P[2]_2 ), .I3(\r_raddr_1P[3]_2 ), .O(n1070)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3900.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3901 (.I0(\r_raddr_1P[0]_2 ), .I1(\r_raddr_1P[1]_2 ), 
            .I2(\r_raddr_1P[2]_2 ), .I3(\r_raddr_1P[3]_2 ), .O(n2421)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3901.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3902 (.I0(\r_raddr_1P[4]_2 ), .I1(n2421), .O(n1075)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3902.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3903 (.I0(\r_raddr_1P[4]_2 ), .I1(n2421), .I2(\r_raddr_1P[5]_2 ), 
            .O(n1080)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3903.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3904 (.I0(\r_raddr_1P[4]_2 ), .I1(\r_raddr_1P[5]_2 ), 
            .O(n2422)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8888 */ ;
    defparam LUT__3904.LUTMASK = 16'h8888;
    EFX_LUT4 LUT__3905 (.I0(n2421), .I1(n2422), .I2(\r_raddr_1P[6]_2 ), 
            .O(n1085)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3905.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3906 (.I0(\r_raddr_1P[6]_2 ), .I1(n2421), .I2(n2422), 
            .I3(\r_raddr_1P[7]_2 ), .O(n1090)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3906.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3907 (.I0(\r_raddr_1P[6]_2 ), .I1(\r_raddr_1P[7]_2 ), 
            .I2(n2421), .I3(n2422), .O(n2423)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3907.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3908 (.I0(\r_raddr_1P[8]_2 ), .I1(n2423), .O(n1095)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3908.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3909 (.I0(\r_raddr_1P[8]_2 ), .I1(n2423), .I2(\r_raddr_1P[9]_2 ), 
            .O(n1100)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3909.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3910 (.I0(\r_raddr_1P[8]_2 ), .I1(\r_raddr_1P[9]_2 ), 
            .I2(n2423), .I3(\r_raddr_1P[10]_2 ), .O(n1105)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7f80 */ ;
    defparam LUT__3910.LUTMASK = 16'h7f80;
    EFX_LUT4 LUT__3911 (.I0(\r_raddr_1P[8]_2 ), .I1(\r_raddr_1P[9]_2 ), 
            .I2(\r_raddr_1P[10]_2 ), .I3(n2423), .O(n2424)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h8000 */ ;
    defparam LUT__3911.LUTMASK = 16'h8000;
    EFX_LUT4 LUT__3912 (.I0(\r_raddr_1P[11]_2 ), .I1(n2424), .O(n1110)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h6666 */ ;
    defparam LUT__3912.LUTMASK = 16'h6666;
    EFX_LUT4 LUT__3913 (.I0(\r_raddr_1P[11]_2 ), .I1(n2424), .I2(\r_raddr_1P[12]_2 ), 
            .O(n1115)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h7878 */ ;
    defparam LUT__3913.LUTMASK = 16'h7878;
    EFX_LUT4 LUT__3914 (.I0(\r_raddr_1P[12]_2 ), .I1(r_rden_1P_2), .O(n1504)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h4444 */ ;
    defparam LUT__3914.LUTMASK = 16'h4444;
    EFX_LUT4 LUT__3915 (.I0(\inst_dly/n29 ), .I1(\inst_dly/n28 ), .I2(\inst_dly/n24 ), 
            .O(\inst_dly/r_rdata_1P[0] )) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hcaca */ ;
    defparam LUT__3915.LUTMASK = 16'hcaca;
    EFX_LUT4 LUT__3916 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[13] ), 
            .O(n2221)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3916.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3917 (.I0(\red_gain[1] ), .I1(\r_mipi_rx_data_1P[12] ), 
            .O(n2223)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3917.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3918 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[39] ), 
            .O(n2278)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3918.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3919 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[38] ), 
            .O(n2281)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3919.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3920 (.I0(\red_gain[0] ), .I1(\r_mipi_rx_data_1P[37] ), 
            .O(n2284)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'hbbbb */ ;
    defparam LUT__3920.LUTMASK = 16'hbbbb;
    EFX_LUT4 LUT__3515 (.I0(\key1_counter[0]_2 ), .I1(\key1_counter[1] ), 
            .I2(\key1_counter[2] ), .I3(\key1_counter[3] ), .O(n2330)) /* verific EFX_ATTRIBUTE_CELL_NAME=EFX_LUT4, LUTMASK=16'h0001 */ ;
    defparam LUT__3515.LUTMASK = 16'h0001;
    
endmodule

//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_237
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_238
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_239
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_240
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_241
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_242
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_243
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_244
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_245
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_246
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_247
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_248
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_249
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_250
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_251
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_252
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_253
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_254
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_255
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_256
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_257
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_258
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_259
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_260
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_261
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_262
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_263
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_264
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_265
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_266
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_267
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_268
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_269
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_270
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_271
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_272
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_273
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_274
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_275
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_276
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_277
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_278
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_279
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_280
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_281
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_282
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_283
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_284
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_285
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_286
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_287
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_288
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_289
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_290
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_291
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_292
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_293
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_294
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_295
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_296
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_297
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_298
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_299
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_300
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_301
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_302
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_303
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_304
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_305
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_306
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_307
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_308
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_309
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_310
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_311
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_312
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_313
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_314
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_315
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_316
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_317
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_318
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_319
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_320
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_321
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_322
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_323
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_324
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_325
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_326
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_327
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_328
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_329
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_330
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_331
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_332
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_333
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_334
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_335
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_336
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_337
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_338
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_339
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_340
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_341
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_342
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_343
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_344
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_345
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_346
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_347
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_348
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_349
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_350
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_351
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_352
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_353
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_354
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_355
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_356
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_357
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_358
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_359
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_360
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_361
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_362
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_363
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_364
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_365
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_366
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_367
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_368
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_369
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_370
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_371
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_372
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_373
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_374
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_375
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_376
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_377
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_378
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_379
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_380
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_381
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_382
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_383
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_384
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_385
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_386
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_387
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_388
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_389
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_390
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_391
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_392
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_393
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_394
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_395
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_396
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_397
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_398
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_399
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_400
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_401
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_402
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_403
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_404
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_405
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_406
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_407
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_408
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_409
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_410
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_411
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_412
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_413
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_414
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_415
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_GBUFCE_c6ffcdc0_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_416
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_417
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_418
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_419
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_420
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_421
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_422
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_423
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_424
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_425
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_426
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_427
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_428
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_FF_c6ffcdc0_429
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_237
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_238
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_239
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_240
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_241
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_242
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_243
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_244
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_245
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_246
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_ADD_c6ffcdc0_247
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_0
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__1_1_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__2_2_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_RAM_5K_c6ffcdc0__1_1_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_1
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_2
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_3
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_4
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_5
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_6
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_7
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_8
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_9
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_10
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_11
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_12
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_13
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_14
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_15
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_16
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_17
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_18
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_19
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_20
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_21
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_22
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_23
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_24
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_25
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_26
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_27
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_28
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_29
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_30
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_31
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_32
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_33
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_34
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_35
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_36
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_37
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_38
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_39
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_40
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_41
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_42
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_43
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_44
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_45
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_46
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_47
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_48
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_49
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_50
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_51
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_52
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_53
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_54
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_55
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_56
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_57
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_58
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_59
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_60
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_61
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_62
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_63
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_64
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_65
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_66
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_67
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_68
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_69
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_70
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_71
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_72
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_73
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_74
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_75
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_76
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_77
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_78
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_79
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_80
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_81
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_82
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_83
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_84
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_85
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_86
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_87
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_88
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_89
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_90
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_91
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_92
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_93
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_94
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_95
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_96
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_97
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_98
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_99
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_100
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_101
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_102
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_103
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_104
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_105
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_106
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_107
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_108
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_109
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_110
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_111
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_112
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_113
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_114
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_115
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_116
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_117
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_118
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_119
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_120
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_121
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_122
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_123
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_124
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_125
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_126
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_127
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_128
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_129
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_130
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_131
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_132
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_133
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_134
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_135
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_136
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_137
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_138
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_139
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_140
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_141
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_142
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_143
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_144
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_145
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_146
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_147
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_148
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_149
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_150
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_151
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_152
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_153
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_154
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_155
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_156
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_157
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_158
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_159
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_160
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_161
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_162
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_163
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_164
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_165
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_166
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_167
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_168
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_169
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_170
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_171
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_172
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_173
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_174
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_175
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_176
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_177
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_178
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_179
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_180
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_181
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_182
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_183
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_184
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_185
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_186
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_187
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_188
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_189
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_190
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_191
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_192
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_193
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_194
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_195
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_196
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_197
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_198
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_199
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_200
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_201
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_202
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_203
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_204
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_205
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_206
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_207
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_208
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_209
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_210
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_211
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_212
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_213
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_214
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_215
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_216
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_217
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_218
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_219
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_220
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_221
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_222
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_223
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_224
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_225
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_226
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_227
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_228
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_229
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_230
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_231
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_232
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_233
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_234
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_235
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_236
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_237
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_238
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_239
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_240
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_241
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_242
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_243
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_244
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_245
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_246
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_247
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_248
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_249
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_250
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_251
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_252
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_253
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_254
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_255
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_256
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_257
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_258
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_259
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_260
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_261
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_262
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_263
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_264
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_265
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_266
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_267
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_268
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_269
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_270
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_271
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_272
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_273
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_274
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_275
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_276
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_277
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_278
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_279
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_280
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_281
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_282
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_283
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_284
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_285
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_286
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_287
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_288
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_289
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_290
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_291
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_292
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_293
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_294
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_295
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_296
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_297
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_298
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_299
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_300
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_301
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_302
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_303
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_304
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_305
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_306
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_307
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_308
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_309
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_310
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_311
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_312
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_313
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_314
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_315
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_316
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_317
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_318
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_319
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_320
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_321
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_322
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_323
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_324
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_325
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_326
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_327
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_328
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_329
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_330
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_331
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_332
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_333
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_334
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_335
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_336
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_337
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_338
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_339
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_340
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_341
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_342
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_343
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_344
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_345
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_346
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_347
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_348
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_349
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_350
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_351
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_352
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_353
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_354
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_355
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_356
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_357
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_358
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_359
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_360
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_361
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_362
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_363
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_364
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_365
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_366
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_367
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_368
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_369
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_370
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_371
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_372
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_373
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_374
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_375
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_376
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_377
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_378
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_379
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_380
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_381
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_382
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_383
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_384
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_385
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_386
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_387
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_388
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_389
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_390
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_391
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_392
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_393
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_394
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_395
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_396
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_397
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_398
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_399
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_400
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_401
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_402
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_403
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_404
// module not written out since it is a black box. 
//


//
// Verific Verilog Description of module EFX_LUT4_c6ffcdc0_405
// module not written out since it is a black box. 
//

